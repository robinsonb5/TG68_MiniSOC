library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity HelloWorld_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1'
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1';
);
end HelloWorld_ROM;

architecture arch of HelloWorld_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))-1) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"ff",
     3 => x"fe",
     4 => x"00",
     5 => x"00",
     6 => x"01",
     7 => x"00",
     8 => x"00",
     9 => x"00",
    10 => x"00",
    11 => x"00",
    12 => x"00",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"00",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"00",
    21 => x"00",
    22 => x"00",
    23 => x"00",
    24 => x"00",
    25 => x"00",
    26 => x"00",
    27 => x"00",
    28 => x"00",
    29 => x"00",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"00",
    34 => x"00",
    35 => x"00",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"00",
    40 => x"00",
    41 => x"00",
    42 => x"00",
    43 => x"00",
    44 => x"00",
    45 => x"00",
    46 => x"00",
    47 => x"00",
    48 => x"00",
    49 => x"00",
    50 => x"00",
    51 => x"00",
    52 => x"00",
    53 => x"00",
    54 => x"00",
    55 => x"00",
    56 => x"00",
    57 => x"00",
    58 => x"00",
    59 => x"00",
    60 => x"00",
    61 => x"00",
    62 => x"00",
    63 => x"00",
    64 => x"00",
    65 => x"00",
    66 => x"00",
    67 => x"00",
    68 => x"00",
    69 => x"00",
    70 => x"00",
    71 => x"00",
    72 => x"00",
    73 => x"00",
    74 => x"00",
    75 => x"00",
    76 => x"00",
    77 => x"00",
    78 => x"00",
    79 => x"00",
    80 => x"00",
    81 => x"00",
    82 => x"00",
    83 => x"00",
    84 => x"00",
    85 => x"00",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"00",
    93 => x"00",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"00",
   127 => x"00",
   128 => x"00",
   129 => x"00",
   130 => x"00",
   131 => x"00",
   132 => x"00",
   133 => x"00",
   134 => x"00",
   135 => x"00",
   136 => x"00",
   137 => x"00",
   138 => x"00",
   139 => x"00",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"00",
   144 => x"00",
   145 => x"00",
   146 => x"00",
   147 => x"00",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"00",
   153 => x"00",
   154 => x"00",
   155 => x"00",
   156 => x"00",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"00",
   161 => x"00",
   162 => x"00",
   163 => x"00",
   164 => x"00",
   165 => x"00",
   166 => x"00",
   167 => x"00",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"00",
   172 => x"00",
   173 => x"00",
   174 => x"00",
   175 => x"00",
   176 => x"00",
   177 => x"00",
   178 => x"00",
   179 => x"00",
   180 => x"00",
   181 => x"00",
   182 => x"00",
   183 => x"00",
   184 => x"00",
   185 => x"00",
   186 => x"00",
   187 => x"00",
   188 => x"00",
   189 => x"00",
   190 => x"00",
   191 => x"00",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"00",
   196 => x"00",
   197 => x"00",
   198 => x"00",
   199 => x"00",
   200 => x"00",
   201 => x"00",
   202 => x"00",
   203 => x"00",
   204 => x"00",
   205 => x"00",
   206 => x"00",
   207 => x"00",
   208 => x"00",
   209 => x"00",
   210 => x"00",
   211 => x"00",
   212 => x"00",
   213 => x"00",
   214 => x"00",
   215 => x"00",
   216 => x"00",
   217 => x"00",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"00",
   224 => x"00",
   225 => x"00",
   226 => x"00",
   227 => x"00",
   228 => x"00",
   229 => x"00",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"00",
   234 => x"00",
   235 => x"00",
   236 => x"00",
   237 => x"00",
   238 => x"00",
   239 => x"00",
   240 => x"00",
   241 => x"00",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"00",
   248 => x"00",
   249 => x"00",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"00",
   256 => x"4f",
   257 => x"f9",
   258 => x"00",
   259 => x"7f",
   260 => x"ff",
   261 => x"fe",
   262 => x"41",
   263 => x"f9",
   264 => x"00",
   265 => x"00",
   266 => x"02",
   267 => x"e0",
   268 => x"20",
   269 => x"3c",
   270 => x"00",
   271 => x"00",
   272 => x"02",
   273 => x"e0",
   274 => x"b1",
   275 => x"c0",
   276 => x"6c",
   277 => x"04",
   278 => x"42",
   279 => x"98",
   280 => x"60",
   281 => x"f8",
   282 => x"41",
   283 => x"fa",
   284 => x"00",
   285 => x"3c",
   286 => x"21",
   287 => x"c8",
   288 => x"00",
   289 => x"64",
   290 => x"41",
   291 => x"fa",
   292 => x"00",
   293 => x"42",
   294 => x"21",
   295 => x"c8",
   296 => x"00",
   297 => x"68",
   298 => x"41",
   299 => x"fa",
   300 => x"00",
   301 => x"48",
   302 => x"21",
   303 => x"c8",
   304 => x"00",
   305 => x"6c",
   306 => x"41",
   307 => x"fa",
   308 => x"00",
   309 => x"4e",
   310 => x"21",
   311 => x"c8",
   312 => x"00",
   313 => x"70",
   314 => x"41",
   315 => x"fa",
   316 => x"00",
   317 => x"54",
   318 => x"21",
   319 => x"c8",
   320 => x"00",
   321 => x"74",
   322 => x"41",
   323 => x"fa",
   324 => x"00",
   325 => x"5a",
   326 => x"21",
   327 => x"c8",
   328 => x"00",
   329 => x"78",
   330 => x"41",
   331 => x"fa",
   332 => x"00",
   333 => x"60",
   334 => x"21",
   335 => x"c8",
   336 => x"00",
   337 => x"7c",
   338 => x"4e",
   339 => x"f9",
   340 => x"00",
   341 => x"00",
   342 => x"02",
   343 => x"70",
   344 => x"48",
   345 => x"e7",
   346 => x"ff",
   347 => x"fe",
   348 => x"48",
   349 => x"7a",
   350 => x"00",
   351 => x"5c",
   352 => x"2f",
   353 => x"3a",
   354 => x"00",
   355 => x"60",
   356 => x"4e",
   357 => x"75",
   358 => x"48",
   359 => x"e7",
   360 => x"ff",
   361 => x"fe",
   362 => x"48",
   363 => x"7a",
   364 => x"00",
   365 => x"4e",
   366 => x"2f",
   367 => x"3a",
   368 => x"00",
   369 => x"56",
   370 => x"4e",
   371 => x"75",
   372 => x"48",
   373 => x"e7",
   374 => x"ff",
   375 => x"fe",
   376 => x"48",
   377 => x"7a",
   378 => x"00",
   379 => x"40",
   380 => x"2f",
   381 => x"3a",
   382 => x"00",
   383 => x"4c",
   384 => x"4e",
   385 => x"75",
   386 => x"48",
   387 => x"e7",
   388 => x"ff",
   389 => x"fe",
   390 => x"48",
   391 => x"7a",
   392 => x"00",
   393 => x"32",
   394 => x"2f",
   395 => x"3a",
   396 => x"00",
   397 => x"42",
   398 => x"4e",
   399 => x"75",
   400 => x"48",
   401 => x"e7",
   402 => x"ff",
   403 => x"fe",
   404 => x"48",
   405 => x"7a",
   406 => x"00",
   407 => x"24",
   408 => x"2f",
   409 => x"3a",
   410 => x"00",
   411 => x"38",
   412 => x"4e",
   413 => x"75",
   414 => x"48",
   415 => x"e7",
   416 => x"ff",
   417 => x"fe",
   418 => x"48",
   419 => x"7a",
   420 => x"00",
   421 => x"16",
   422 => x"2f",
   423 => x"3a",
   424 => x"00",
   425 => x"2e",
   426 => x"4e",
   427 => x"75",
   428 => x"48",
   429 => x"e7",
   430 => x"ff",
   431 => x"fe",
   432 => x"48",
   433 => x"7a",
   434 => x"00",
   435 => x"08",
   436 => x"2f",
   437 => x"3a",
   438 => x"00",
   439 => x"24",
   440 => x"4e",
   441 => x"75",
   442 => x"4c",
   443 => x"df",
   444 => x"7f",
   445 => x"ff",
   446 => x"4e",
   447 => x"73",
   448 => x"4e",
   449 => x"75",
   450 => x"00",
   451 => x"00",
   452 => x"01",
   453 => x"c0",
   454 => x"00",
   455 => x"00",
   456 => x"01",
   457 => x"c0",
   458 => x"00",
   459 => x"00",
   460 => x"01",
   461 => x"c0",
   462 => x"00",
   463 => x"00",
   464 => x"01",
   465 => x"c0",
   466 => x"00",
   467 => x"00",
   468 => x"01",
   469 => x"c0",
   470 => x"00",
   471 => x"00",
   472 => x"01",
   473 => x"c0",
   474 => x"00",
   475 => x"00",
   476 => x"01",
   477 => x"c0",
   478 => x"46",
   479 => x"fc",
   480 => x"20",
   481 => x"00",
   482 => x"4e",
   483 => x"75",
   484 => x"46",
   485 => x"fc",
   486 => x"27",
   487 => x"00",
   488 => x"4e",
   489 => x"75",
   490 => x"00",
   491 => x"00",
   492 => x"00",
   493 => x"00",
   494 => x"00",
   495 => x"00",
   496 => x"cf",
   497 => x"00",
   498 => x"00",
   499 => x"00",
   500 => x"00",
   501 => x"00",
   502 => x"00",
   503 => x"00",
   504 => x"8c",
   505 => x"ff",
   506 => x"f0",
   507 => x"00",
   508 => x"00",
   509 => x"00",
   510 => x"00",
   511 => x"00",
   512 => x"08",
   513 => x"cc",
   514 => x"ff",
   515 => x"f0",
   516 => x"00",
   517 => x"00",
   518 => x"00",
   519 => x"00",
   520 => x"08",
   521 => x"cc",
   522 => x"cc",
   523 => x"ff",
   524 => x"ff",
   525 => x"00",
   526 => x"00",
   527 => x"00",
   528 => x"08",
   529 => x"8c",
   530 => x"cc",
   531 => x"cc",
   532 => x"cf",
   533 => x"ff",
   534 => x"00",
   535 => x"00",
   536 => x"00",
   537 => x"8c",
   538 => x"cc",
   539 => x"cc",
   540 => x"cc",
   541 => x"c8",
   542 => x"00",
   543 => x"00",
   544 => x"00",
   545 => x"88",
   546 => x"cc",
   547 => x"cc",
   548 => x"cc",
   549 => x"80",
   550 => x"00",
   551 => x"00",
   552 => x"00",
   553 => x"08",
   554 => x"cc",
   555 => x"cc",
   556 => x"cf",
   557 => x"00",
   558 => x"00",
   559 => x"00",
   560 => x"00",
   561 => x"08",
   562 => x"cc",
   563 => x"cc",
   564 => x"cc",
   565 => x"f0",
   566 => x"00",
   567 => x"00",
   568 => x"00",
   569 => x"08",
   570 => x"8c",
   571 => x"c8",
   572 => x"cc",
   573 => x"cf",
   574 => x"00",
   575 => x"00",
   576 => x"00",
   577 => x"00",
   578 => x"8c",
   579 => x"80",
   580 => x"8c",
   581 => x"cc",
   582 => x"f0",
   583 => x"00",
   584 => x"00",
   585 => x"00",
   586 => x"88",
   587 => x"00",
   588 => x"08",
   589 => x"cc",
   590 => x"cf",
   591 => x"00",
   592 => x"00",
   593 => x"00",
   594 => x"00",
   595 => x"00",
   596 => x"00",
   597 => x"8c",
   598 => x"cc",
   599 => x"f0",
   600 => x"00",
   601 => x"00",
   602 => x"00",
   603 => x"00",
   604 => x"00",
   605 => x"08",
   606 => x"cc",
   607 => x"c8",
   608 => x"00",
   609 => x"00",
   610 => x"00",
   611 => x"00",
   612 => x"00",
   613 => x"00",
   614 => x"8c",
   615 => x"80",
   616 => x"00",
   617 => x"00",
   618 => x"00",
   619 => x"00",
   620 => x"00",
   621 => x"00",
   622 => x"08",
   623 => x"00",
   624 => x"4e",
   625 => x"56",
   626 => x"00",
   627 => x"00",
   628 => x"48",
   629 => x"79",
   630 => x"00",
   631 => x"00",
   632 => x"02",
   633 => x"ce",
   634 => x"4e",
   635 => x"b9",
   636 => x"00",
   637 => x"00",
   638 => x"02",
   639 => x"a2",
   640 => x"42",
   641 => x"80",
   642 => x"4e",
   643 => x"5e",
   644 => x"4e",
   645 => x"75",
   646 => x"00",
   647 => x"00",
   648 => x"4e",
   649 => x"56",
   650 => x"00",
   651 => x"00",
   652 => x"20",
   653 => x"2e",
   654 => x"00",
   655 => x"08",
   656 => x"22",
   657 => x"38",
   658 => x"ff",
   659 => x"c0",
   660 => x"08",
   661 => x"01",
   662 => x"00",
   663 => x"08",
   664 => x"67",
   665 => x"f6",
   666 => x"21",
   667 => x"c0",
   668 => x"ff",
   669 => x"c0",
   670 => x"4e",
   671 => x"5e",
   672 => x"4e",
   673 => x"75",
   674 => x"4e",
   675 => x"56",
   676 => x"00",
   677 => x"00",
   678 => x"48",
   679 => x"e7",
   680 => x"20",
   681 => x"30",
   682 => x"24",
   683 => x"6e",
   684 => x"00",
   685 => x"08",
   686 => x"47",
   687 => x"fa",
   688 => x"ff",
   689 => x"d8",
   690 => x"60",
   691 => x"0a",
   692 => x"49",
   693 => x"c0",
   694 => x"2f",
   695 => x"00",
   696 => x"4e",
   697 => x"93",
   698 => x"52",
   699 => x"82",
   700 => x"58",
   701 => x"8f",
   702 => x"10",
   703 => x"1a",
   704 => x"66",
   705 => x"f2",
   706 => x"20",
   707 => x"02",
   708 => x"4c",
   709 => x"ee",
   710 => x"0c",
   711 => x"04",
   712 => x"ff",
   713 => x"f4",
   714 => x"4e",
   715 => x"5e",
   716 => x"4e",
   717 => x"75",
   718 => x"48",
   719 => x"65",
   720 => x"6c",
   721 => x"6c",
   722 => x"6f",
   723 => x"2c",
   724 => x"20",
   725 => x"77",
   726 => x"6f",
   727 => x"72",
   728 => x"6c",
   729 => x"64",
   730 => x"21",
   731 => x"0a",
   732 => x"00",
   733 => x"00",
   734 => x"00",
   735 => x"00",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we = '0' and lds='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we = '0' and uds='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


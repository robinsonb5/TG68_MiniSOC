library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"41",
    49 => x"fa",
    50 => x"00",
    51 => x"74",
    52 => x"61",
    53 => x"00",
    54 => x"02",
    55 => x"d8",
    56 => x"33",
    57 => x"fc",
    58 => x"0f",
    59 => x"00",
    60 => x"81",
    61 => x"00",
    62 => x"00",
    63 => x"06",
    64 => x"2e",
    65 => x"3c",
    66 => x"00",
    67 => x"00",
    68 => x"07",
    69 => x"ff",
    70 => x"41",
    71 => x"f9",
    72 => x"80",
    73 => x"00",
    74 => x"08",
    75 => x"00",
    76 => x"10",
    77 => x"fc",
    78 => x"00",
    79 => x"20",
    80 => x"51",
    81 => x"cf",
    82 => x"ff",
    83 => x"fa",
    84 => x"23",
    85 => x"fc",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"7f",
    92 => x"00",
    93 => x"52",
    94 => x"41",
    95 => x"fa",
    96 => x"00",
    97 => x"46",
    98 => x"61",
    99 => x"00",
   100 => x"06",
   101 => x"ba",
   102 => x"61",
   103 => x"00",
   104 => x"0a",
   105 => x"ec",
   106 => x"4a",
   107 => x"80",
   108 => x"67",
   109 => x"0a",
   110 => x"41",
   111 => x"fa",
   112 => x"00",
   113 => x"6a",
   114 => x"61",
   115 => x"00",
   116 => x"06",
   117 => x"aa",
   118 => x"60",
   119 => x"fe",
   120 => x"41",
   121 => x"fa",
   122 => x"00",
   123 => x"49",
   124 => x"61",
   125 => x"00",
   126 => x"06",
   127 => x"a0",
   128 => x"61",
   129 => x"00",
   130 => x"02",
   131 => x"ac",
   132 => x"4b",
   133 => x"f9",
   134 => x"80",
   135 => x"00",
   136 => x"08",
   137 => x"00",
   138 => x"33",
   139 => x"fc",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"7f",
   144 => x"00",
   145 => x"0c",
   146 => x"30",
   147 => x"39",
   148 => x"81",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"08",
   153 => x"00",
   154 => x"00",
   155 => x"09",
   156 => x"67",
   157 => x"f4",
   158 => x"3a",
   159 => x"c0",
   160 => x"61",
   161 => x"00",
   162 => x"00",
   163 => x"80",
   164 => x"60",
   165 => x"ec",
   166 => x"43",
   167 => x"6f",
   168 => x"6e",
   169 => x"64",
   170 => x"75",
   171 => x"63",
   172 => x"74",
   173 => x"69",
   174 => x"6e",
   175 => x"67",
   176 => x"20",
   177 => x"73",
   178 => x"61",
   179 => x"6e",
   180 => x"69",
   181 => x"74",
   182 => x"79",
   183 => x"20",
   184 => x"63",
   185 => x"68",
   186 => x"65",
   187 => x"63",
   188 => x"6b",
   189 => x"2e",
   190 => x"2e",
   191 => x"2e",
   192 => x"0d",
   193 => x"0a",
   194 => x"00",
   195 => x"53",
   196 => x"61",
   197 => x"6e",
   198 => x"69",
   199 => x"74",
   200 => x"79",
   201 => x"20",
   202 => x"63",
   203 => x"68",
   204 => x"65",
   205 => x"63",
   206 => x"6b",
   207 => x"20",
   208 => x"70",
   209 => x"61",
   210 => x"73",
   211 => x"73",
   212 => x"65",
   213 => x"64",
   214 => x"2e",
   215 => x"0d",
   216 => x"0a",
   217 => x"00",
   218 => x"53",
   219 => x"61",
   220 => x"6e",
   221 => x"69",
   222 => x"74",
   223 => x"79",
   224 => x"20",
   225 => x"63",
   226 => x"68",
   227 => x"65",
   228 => x"63",
   229 => x"6b",
   230 => x"20",
   231 => x"66",
   232 => x"61",
   233 => x"69",
   234 => x"6c",
   235 => x"65",
   236 => x"64",
   237 => x"2e",
   238 => x"0d",
   239 => x"0a",
   240 => x"00",
   241 => x"00",
   242 => x"c0",
   243 => x"bc",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"df",
   248 => x"90",
   249 => x"3c",
   250 => x"00",
   251 => x"37",
   252 => x"6a",
   253 => x"04",
   254 => x"d0",
   255 => x"3c",
   256 => x"00",
   257 => x"27",
   258 => x"e9",
   259 => x"8e",
   260 => x"8c",
   261 => x"00",
   262 => x"20",
   263 => x"86",
   264 => x"4e",
   265 => x"75",
   266 => x"c0",
   267 => x"bc",
   268 => x"00",
   269 => x"00",
   270 => x"00",
   271 => x"df",
   272 => x"90",
   273 => x"3c",
   274 => x"00",
   275 => x"37",
   276 => x"6a",
   277 => x"04",
   278 => x"d0",
   279 => x"3c",
   280 => x"00",
   281 => x"27",
   282 => x"e9",
   283 => x"0f",
   284 => x"8e",
   285 => x"00",
   286 => x"10",
   287 => x"87",
   288 => x"4e",
   289 => x"75",
   290 => x"52",
   291 => x"79",
   292 => x"00",
   293 => x"7f",
   294 => x"00",
   295 => x"0c",
   296 => x"b0",
   297 => x"3c",
   298 => x"00",
   299 => x"53",
   300 => x"66",
   301 => x"2a",
   302 => x"33",
   303 => x"fc",
   304 => x"ff",
   305 => x"ff",
   306 => x"81",
   307 => x"00",
   308 => x"00",
   309 => x"06",
   310 => x"72",
   311 => x"00",
   312 => x"2e",
   313 => x"01",
   314 => x"2c",
   315 => x"01",
   316 => x"33",
   317 => x"c1",
   318 => x"00",
   319 => x"7f",
   320 => x"00",
   321 => x"0c",
   322 => x"23",
   323 => x"c1",
   324 => x"00",
   325 => x"7f",
   326 => x"00",
   327 => x"08",
   328 => x"23",
   329 => x"c1",
   330 => x"00",
   331 => x"7f",
   332 => x"00",
   333 => x"04",
   334 => x"23",
   335 => x"c1",
   336 => x"00",
   337 => x"7f",
   338 => x"00",
   339 => x"10",
   340 => x"60",
   341 => x"00",
   342 => x"01",
   343 => x"72",
   344 => x"2c",
   345 => x"39",
   346 => x"00",
   347 => x"7f",
   348 => x"00",
   349 => x"20",
   350 => x"2e",
   351 => x"39",
   352 => x"00",
   353 => x"7f",
   354 => x"00",
   355 => x"1c",
   356 => x"0c",
   357 => x"79",
   358 => x"00",
   359 => x"01",
   360 => x"00",
   361 => x"7f",
   362 => x"00",
   363 => x"0c",
   364 => x"66",
   365 => x"34",
   366 => x"33",
   367 => x"fc",
   368 => x"f0",
   369 => x"00",
   370 => x"81",
   371 => x"00",
   372 => x"00",
   373 => x"06",
   374 => x"41",
   375 => x"f9",
   376 => x"00",
   377 => x"7f",
   378 => x"00",
   379 => x"13",
   380 => x"61",
   381 => x"8c",
   382 => x"22",
   383 => x"39",
   384 => x"00",
   385 => x"7f",
   386 => x"00",
   387 => x"10",
   388 => x"b2",
   389 => x"bc",
   390 => x"00",
   391 => x"00",
   392 => x"00",
   393 => x"03",
   394 => x"6f",
   395 => x"08",
   396 => x"72",
   397 => x"0a",
   398 => x"92",
   399 => x"b9",
   400 => x"00",
   401 => x"7f",
   402 => x"00",
   403 => x"10",
   404 => x"52",
   405 => x"81",
   406 => x"e3",
   407 => x"89",
   408 => x"23",
   409 => x"c1",
   410 => x"00",
   411 => x"7f",
   412 => x"00",
   413 => x"14",
   414 => x"60",
   415 => x"00",
   416 => x"01",
   417 => x"28",
   418 => x"33",
   419 => x"f9",
   420 => x"00",
   421 => x"7f",
   422 => x"00",
   423 => x"12",
   424 => x"81",
   425 => x"00",
   426 => x"00",
   427 => x"06",
   428 => x"4a",
   429 => x"b9",
   430 => x"00",
   431 => x"7f",
   432 => x"00",
   433 => x"10",
   434 => x"67",
   435 => x"00",
   436 => x"01",
   437 => x"14",
   438 => x"0c",
   439 => x"b9",
   440 => x"00",
   441 => x"00",
   442 => x"00",
   443 => x"09",
   444 => x"00",
   445 => x"7f",
   446 => x"00",
   447 => x"10",
   448 => x"6e",
   449 => x"00",
   450 => x"00",
   451 => x"c0",
   452 => x"0c",
   453 => x"79",
   454 => x"00",
   455 => x"03",
   456 => x"00",
   457 => x"7f",
   458 => x"00",
   459 => x"0c",
   460 => x"6e",
   461 => x"16",
   462 => x"33",
   463 => x"fc",
   464 => x"0f",
   465 => x"00",
   466 => x"81",
   467 => x"00",
   468 => x"00",
   469 => x"06",
   470 => x"41",
   471 => x"f9",
   472 => x"00",
   473 => x"7f",
   474 => x"00",
   475 => x"07",
   476 => x"61",
   477 => x"00",
   478 => x"ff",
   479 => x"2c",
   480 => x"60",
   481 => x"00",
   482 => x"00",
   483 => x"e6",
   484 => x"22",
   485 => x"39",
   486 => x"00",
   487 => x"7f",
   488 => x"00",
   489 => x"14",
   490 => x"56",
   491 => x"41",
   492 => x"34",
   493 => x"39",
   494 => x"00",
   495 => x"7f",
   496 => x"00",
   497 => x"0c",
   498 => x"b4",
   499 => x"41",
   500 => x"6e",
   501 => x"20",
   502 => x"41",
   503 => x"f9",
   504 => x"00",
   505 => x"7f",
   506 => x"00",
   507 => x"08",
   508 => x"61",
   509 => x"00",
   510 => x"fe",
   511 => x"f4",
   512 => x"33",
   513 => x"f9",
   514 => x"00",
   515 => x"7f",
   516 => x"00",
   517 => x"0a",
   518 => x"81",
   519 => x"00",
   520 => x"00",
   521 => x"06",
   522 => x"33",
   523 => x"fc",
   524 => x"00",
   525 => x"01",
   526 => x"00",
   527 => x"7f",
   528 => x"00",
   529 => x"18",
   530 => x"60",
   531 => x"00",
   532 => x"00",
   533 => x"b4",
   534 => x"0c",
   535 => x"b9",
   536 => x"00",
   537 => x"00",
   538 => x"00",
   539 => x"03",
   540 => x"00",
   541 => x"7f",
   542 => x"00",
   543 => x"10",
   544 => x"6e",
   545 => x"60",
   546 => x"33",
   547 => x"fc",
   548 => x"00",
   549 => x"0f",
   550 => x"81",
   551 => x"00",
   552 => x"00",
   553 => x"06",
   554 => x"22",
   555 => x"39",
   556 => x"00",
   557 => x"7f",
   558 => x"00",
   559 => x"04",
   560 => x"e3",
   561 => x"89",
   562 => x"52",
   563 => x"81",
   564 => x"34",
   565 => x"39",
   566 => x"00",
   567 => x"7f",
   568 => x"00",
   569 => x"0c",
   570 => x"b4",
   571 => x"41",
   572 => x"6e",
   573 => x"2a",
   574 => x"20",
   575 => x"79",
   576 => x"00",
   577 => x"7f",
   578 => x"00",
   579 => x"08",
   580 => x"61",
   581 => x"00",
   582 => x"fe",
   583 => x"c4",
   584 => x"32",
   585 => x"39",
   586 => x"00",
   587 => x"7f",
   588 => x"00",
   589 => x"18",
   590 => x"53",
   591 => x"79",
   592 => x"00",
   593 => x"7f",
   594 => x"00",
   595 => x"18",
   596 => x"53",
   597 => x"41",
   598 => x"6a",
   599 => x"70",
   600 => x"52",
   601 => x"b9",
   602 => x"00",
   603 => x"7f",
   604 => x"00",
   605 => x"08",
   606 => x"33",
   607 => x"fc",
   608 => x"00",
   609 => x"01",
   610 => x"00",
   611 => x"7f",
   612 => x"00",
   613 => x"18",
   614 => x"60",
   615 => x"60",
   616 => x"30",
   617 => x"39",
   618 => x"00",
   619 => x"7f",
   620 => x"00",
   621 => x"18",
   622 => x"52",
   623 => x"40",
   624 => x"c0",
   625 => x"7c",
   626 => x"00",
   627 => x"01",
   628 => x"67",
   629 => x"52",
   630 => x"20",
   631 => x"79",
   632 => x"00",
   633 => x"7f",
   634 => x"00",
   635 => x"08",
   636 => x"e5",
   637 => x"88",
   638 => x"e1",
   639 => x"2f",
   640 => x"10",
   641 => x"87",
   642 => x"33",
   643 => x"fc",
   644 => x"f0",
   645 => x"f0",
   646 => x"81",
   647 => x"00",
   648 => x"00",
   649 => x"06",
   650 => x"0c",
   651 => x"b9",
   652 => x"00",
   653 => x"00",
   654 => x"00",
   655 => x"07",
   656 => x"00",
   657 => x"7f",
   658 => x"00",
   659 => x"10",
   660 => x"6d",
   661 => x"32",
   662 => x"33",
   663 => x"fc",
   664 => x"f0",
   665 => x"0f",
   666 => x"81",
   667 => x"00",
   668 => x"00",
   669 => x"06",
   670 => x"0c",
   671 => x"b9",
   672 => x"00",
   673 => x"00",
   674 => x"00",
   675 => x"09",
   676 => x"00",
   677 => x"7f",
   678 => x"00",
   679 => x"10",
   680 => x"6e",
   681 => x"1e",
   682 => x"33",
   683 => x"fc",
   684 => x"ff",
   685 => x"f0",
   686 => x"81",
   687 => x"00",
   688 => x"00",
   689 => x"06",
   690 => x"41",
   691 => x"fa",
   692 => x"00",
   693 => x"22",
   694 => x"61",
   695 => x"56",
   696 => x"2e",
   697 => x"b9",
   698 => x"00",
   699 => x"7f",
   700 => x"00",
   701 => x"08",
   702 => x"08",
   703 => x"b9",
   704 => x"00",
   705 => x"00",
   706 => x"81",
   707 => x"00",
   708 => x"00",
   709 => x"04",
   710 => x"4e",
   711 => x"75",
   712 => x"23",
   713 => x"c6",
   714 => x"00",
   715 => x"7f",
   716 => x"00",
   717 => x"20",
   718 => x"23",
   719 => x"c7",
   720 => x"00",
   721 => x"7f",
   722 => x"00",
   723 => x"1c",
   724 => x"4e",
   725 => x"75",
   726 => x"46",
   727 => x"69",
   728 => x"72",
   729 => x"6d",
   730 => x"77",
   731 => x"61",
   732 => x"72",
   733 => x"65",
   734 => x"20",
   735 => x"72",
   736 => x"65",
   737 => x"63",
   738 => x"65",
   739 => x"69",
   740 => x"76",
   741 => x"65",
   742 => x"64",
   743 => x"20",
   744 => x"2d",
   745 => x"20",
   746 => x"6c",
   747 => x"61",
   748 => x"75",
   749 => x"6e",
   750 => x"63",
   751 => x"68",
   752 => x"69",
   753 => x"6e",
   754 => x"67",
   755 => x"0d",
   756 => x"0a",
   757 => x"00",
   758 => x"48",
   759 => x"40",
   760 => x"30",
   761 => x"39",
   762 => x"81",
   763 => x"00",
   764 => x"00",
   765 => x"00",
   766 => x"08",
   767 => x"00",
   768 => x"00",
   769 => x"08",
   770 => x"67",
   771 => x"f4",
   772 => x"48",
   773 => x"40",
   774 => x"33",
   775 => x"c0",
   776 => x"81",
   777 => x"00",
   778 => x"00",
   779 => x"00",
   780 => x"4e",
   781 => x"75",
   782 => x"2f",
   783 => x"00",
   784 => x"70",
   785 => x"00",
   786 => x"30",
   787 => x"39",
   788 => x"81",
   789 => x"00",
   790 => x"00",
   791 => x"00",
   792 => x"08",
   793 => x"00",
   794 => x"00",
   795 => x"08",
   796 => x"67",
   797 => x"f4",
   798 => x"10",
   799 => x"18",
   800 => x"67",
   801 => x"08",
   802 => x"33",
   803 => x"c0",
   804 => x"81",
   805 => x"00",
   806 => x"00",
   807 => x"00",
   808 => x"60",
   809 => x"e8",
   810 => x"20",
   811 => x"1f",
   812 => x"4e",
   813 => x"75",
   814 => x"33",
   815 => x"fc",
   816 => x"00",
   817 => x"01",
   818 => x"81",
   819 => x"00",
   820 => x"00",
   821 => x"06",
   822 => x"41",
   823 => x"fa",
   824 => x"01",
   825 => x"fa",
   826 => x"61",
   827 => x"00",
   828 => x"03",
   829 => x"e2",
   830 => x"61",
   831 => x"00",
   832 => x"02",
   833 => x"60",
   834 => x"66",
   835 => x"5c",
   836 => x"33",
   837 => x"fc",
   838 => x"00",
   839 => x"02",
   840 => x"81",
   841 => x"00",
   842 => x"00",
   843 => x"06",
   844 => x"33",
   845 => x"fc",
   846 => x"00",
   847 => x"40",
   848 => x"00",
   849 => x"7f",
   850 => x"00",
   851 => x"26",
   852 => x"61",
   853 => x"00",
   854 => x"04",
   855 => x"8a",
   856 => x"67",
   857 => x"0c",
   858 => x"42",
   859 => x"79",
   860 => x"00",
   861 => x"7f",
   862 => x"00",
   863 => x"26",
   864 => x"61",
   865 => x"00",
   866 => x"04",
   867 => x"7e",
   868 => x"66",
   869 => x"28",
   870 => x"33",
   871 => x"fc",
   872 => x"00",
   873 => x"03",
   874 => x"81",
   875 => x"00",
   876 => x"00",
   877 => x"06",
   878 => x"61",
   879 => x"00",
   880 => x"05",
   881 => x"f8",
   882 => x"43",
   883 => x"fa",
   884 => x"00",
   885 => x"57",
   886 => x"61",
   887 => x"00",
   888 => x"06",
   889 => x"48",
   890 => x"67",
   891 => x"12",
   892 => x"41",
   893 => x"fa",
   894 => x"00",
   895 => x"47",
   896 => x"61",
   897 => x"00",
   898 => x"03",
   899 => x"9c",
   900 => x"30",
   901 => x"7c",
   902 => x"20",
   903 => x"00",
   904 => x"61",
   905 => x"00",
   906 => x"04",
   907 => x"02",
   908 => x"4e",
   909 => x"75",
   910 => x"33",
   911 => x"fc",
   912 => x"f0",
   913 => x"03",
   914 => x"81",
   915 => x"00",
   916 => x"00",
   917 => x"06",
   918 => x"41",
   919 => x"fa",
   920 => x"00",
   921 => x"29",
   922 => x"61",
   923 => x"00",
   924 => x"03",
   925 => x"82",
   926 => x"4e",
   927 => x"75",
   928 => x"33",
   929 => x"fc",
   930 => x"f0",
   931 => x"02",
   932 => x"81",
   933 => x"00",
   934 => x"00",
   935 => x"06",
   936 => x"41",
   937 => x"fa",
   938 => x"00",
   939 => x"08",
   940 => x"61",
   941 => x"00",
   942 => x"03",
   943 => x"70",
   944 => x"4e",
   945 => x"75",
   946 => x"53",
   947 => x"44",
   948 => x"20",
   949 => x"69",
   950 => x"6e",
   951 => x"69",
   952 => x"74",
   953 => x"20",
   954 => x"66",
   955 => x"61",
   956 => x"69",
   957 => x"6c",
   958 => x"65",
   959 => x"64",
   960 => x"00",
   961 => x"6e",
   962 => x"6f",
   963 => x"74",
   964 => x"20",
   965 => x"66",
   966 => x"6f",
   967 => x"75",
   968 => x"6e",
   969 => x"64",
   970 => x"20",
   971 => x"42",
   972 => x"4f",
   973 => x"4f",
   974 => x"54",
   975 => x"20",
   976 => x"20",
   977 => x"20",
   978 => x"20",
   979 => x"53",
   980 => x"52",
   981 => x"45",
   982 => x"00",
   983 => x"00",
   984 => x"33",
   985 => x"fc",
   986 => x"01",
   987 => x"00",
   988 => x"81",
   989 => x"00",
   990 => x"00",
   991 => x"06",
   992 => x"41",
   993 => x"f9",
   994 => x"00",
   995 => x"7f",
   996 => x"00",
   997 => x"56",
   998 => x"61",
   999 => x"00",
  1000 => x"00",
  1001 => x"c4",
  1002 => x"66",
  1003 => x"68",
  1004 => x"33",
  1005 => x"fc",
  1006 => x"01",
  1007 => x"01",
  1008 => x"81",
  1009 => x"00",
  1010 => x"00",
  1011 => x"06",
  1012 => x"32",
  1013 => x"3c",
  1014 => x"4e",
  1015 => x"20",
  1016 => x"53",
  1017 => x"41",
  1018 => x"67",
  1019 => x"44",
  1020 => x"33",
  1021 => x"fc",
  1022 => x"01",
  1023 => x"02",
  1024 => x"81",
  1025 => x"00",
  1026 => x"00",
  1027 => x"06",
  1028 => x"33",
  1029 => x"7c",
  1030 => x"00",
  1031 => x"ff",
  1032 => x"00",
  1033 => x"24",
  1034 => x"30",
  1035 => x"29",
  1036 => x"00",
  1037 => x"24",
  1038 => x"b0",
  1039 => x"3c",
  1040 => x"00",
  1041 => x"fe",
  1042 => x"66",
  1043 => x"e4",
  1044 => x"30",
  1045 => x"29",
  1046 => x"01",
  1047 => x"00",
  1048 => x"32",
  1049 => x"3c",
  1050 => x"00",
  1051 => x"7f",
  1052 => x"20",
  1053 => x"29",
  1054 => x"01",
  1055 => x"00",
  1056 => x"20",
  1057 => x"c0",
  1058 => x"51",
  1059 => x"c9",
  1060 => x"ff",
  1061 => x"f8",
  1062 => x"30",
  1063 => x"29",
  1064 => x"00",
  1065 => x"24",
  1066 => x"33",
  1067 => x"7c",
  1068 => x"00",
  1069 => x"00",
  1070 => x"00",
  1071 => x"22",
  1072 => x"33",
  1073 => x"fc",
  1074 => x"01",
  1075 => x"03",
  1076 => x"81",
  1077 => x"00",
  1078 => x"00",
  1079 => x"06",
  1080 => x"41",
  1081 => x"e8",
  1082 => x"fe",
  1083 => x"00",
  1084 => x"70",
  1085 => x"00",
  1086 => x"4e",
  1087 => x"75",
  1088 => x"33",
  1089 => x"fc",
  1090 => x"f1",
  1091 => x"02",
  1092 => x"81",
  1093 => x"00",
  1094 => x"00",
  1095 => x"06",
  1096 => x"41",
  1097 => x"fa",
  1098 => x"01",
  1099 => x"38",
  1100 => x"61",
  1101 => x"00",
  1102 => x"02",
  1103 => x"d0",
  1104 => x"70",
  1105 => x"fe",
  1106 => x"4e",
  1107 => x"75",
  1108 => x"33",
  1109 => x"fc",
  1110 => x"f1",
  1111 => x"03",
  1112 => x"81",
  1113 => x"00",
  1114 => x"00",
  1115 => x"06",
  1116 => x"41",
  1117 => x"fa",
  1118 => x"01",
  1119 => x"0c",
  1120 => x"61",
  1121 => x"00",
  1122 => x"02",
  1123 => x"bc",
  1124 => x"70",
  1125 => x"ff",
  1126 => x"4e",
  1127 => x"75",
  1128 => x"22",
  1129 => x"3c",
  1130 => x"00",
  1131 => x"95",
  1132 => x"00",
  1133 => x"40",
  1134 => x"70",
  1135 => x"00",
  1136 => x"60",
  1137 => x"40",
  1138 => x"22",
  1139 => x"3c",
  1140 => x"00",
  1141 => x"ff",
  1142 => x"00",
  1143 => x"41",
  1144 => x"70",
  1145 => x"00",
  1146 => x"60",
  1147 => x"36",
  1148 => x"22",
  1149 => x"3c",
  1150 => x"00",
  1151 => x"87",
  1152 => x"00",
  1153 => x"48",
  1154 => x"20",
  1155 => x"3c",
  1156 => x"00",
  1157 => x"00",
  1158 => x"01",
  1159 => x"aa",
  1160 => x"60",
  1161 => x"28",
  1162 => x"22",
  1163 => x"3c",
  1164 => x"00",
  1165 => x"87",
  1166 => x"00",
  1167 => x"69",
  1168 => x"20",
  1169 => x"3c",
  1170 => x"40",
  1171 => x"00",
  1172 => x"00",
  1173 => x"00",
  1174 => x"60",
  1175 => x"1a",
  1176 => x"22",
  1177 => x"3c",
  1178 => x"00",
  1179 => x"ff",
  1180 => x"00",
  1181 => x"77",
  1182 => x"70",
  1183 => x"00",
  1184 => x"60",
  1185 => x"10",
  1186 => x"22",
  1187 => x"3c",
  1188 => x"00",
  1189 => x"ff",
  1190 => x"00",
  1191 => x"7a",
  1192 => x"70",
  1193 => x"00",
  1194 => x"60",
  1195 => x"06",
  1196 => x"22",
  1197 => x"3c",
  1198 => x"00",
  1199 => x"ff",
  1200 => x"00",
  1201 => x"51",
  1202 => x"43",
  1203 => x"f9",
  1204 => x"81",
  1205 => x"00",
  1206 => x"00",
  1207 => x"00",
  1208 => x"33",
  1209 => x"7c",
  1210 => x"00",
  1211 => x"ff",
  1212 => x"00",
  1213 => x"24",
  1214 => x"3f",
  1215 => x"69",
  1216 => x"00",
  1217 => x"24",
  1218 => x"ff",
  1219 => x"fe",
  1220 => x"33",
  1221 => x"7c",
  1222 => x"00",
  1223 => x"01",
  1224 => x"00",
  1225 => x"22",
  1226 => x"33",
  1227 => x"7c",
  1228 => x"00",
  1229 => x"ff",
  1230 => x"00",
  1231 => x"24",
  1232 => x"33",
  1233 => x"41",
  1234 => x"00",
  1235 => x"24",
  1236 => x"48",
  1237 => x"41",
  1238 => x"4a",
  1239 => x"79",
  1240 => x"00",
  1241 => x"7f",
  1242 => x"00",
  1243 => x"24",
  1244 => x"67",
  1245 => x"16",
  1246 => x"e1",
  1247 => x"98",
  1248 => x"33",
  1249 => x"40",
  1250 => x"00",
  1251 => x"24",
  1252 => x"e1",
  1253 => x"98",
  1254 => x"33",
  1255 => x"40",
  1256 => x"00",
  1257 => x"24",
  1258 => x"e1",
  1259 => x"98",
  1260 => x"33",
  1261 => x"40",
  1262 => x"00",
  1263 => x"24",
  1264 => x"e1",
  1265 => x"98",
  1266 => x"60",
  1267 => x"18",
  1268 => x"d0",
  1269 => x"80",
  1270 => x"48",
  1271 => x"40",
  1272 => x"33",
  1273 => x"40",
  1274 => x"00",
  1275 => x"24",
  1276 => x"48",
  1277 => x"40",
  1278 => x"e1",
  1279 => x"58",
  1280 => x"33",
  1281 => x"40",
  1282 => x"00",
  1283 => x"24",
  1284 => x"e1",
  1285 => x"58",
  1286 => x"33",
  1287 => x"40",
  1288 => x"00",
  1289 => x"24",
  1290 => x"70",
  1291 => x"00",
  1292 => x"33",
  1293 => x"40",
  1294 => x"00",
  1295 => x"24",
  1296 => x"33",
  1297 => x"41",
  1298 => x"00",
  1299 => x"24",
  1300 => x"22",
  1301 => x"3c",
  1302 => x"00",
  1303 => x"00",
  1304 => x"01",
  1305 => x"90",
  1306 => x"53",
  1307 => x"81",
  1308 => x"67",
  1309 => x"10",
  1310 => x"33",
  1311 => x"7c",
  1312 => x"00",
  1313 => x"ff",
  1314 => x"00",
  1315 => x"24",
  1316 => x"30",
  1317 => x"29",
  1318 => x"00",
  1319 => x"24",
  1320 => x"b0",
  1321 => x"3c",
  1322 => x"00",
  1323 => x"ff",
  1324 => x"67",
  1325 => x"ec",
  1326 => x"80",
  1327 => x"00",
  1328 => x"4e",
  1329 => x"75",
  1330 => x"53",
  1331 => x"74",
  1332 => x"61",
  1333 => x"72",
  1334 => x"74",
  1335 => x"20",
  1336 => x"49",
  1337 => x"6e",
  1338 => x"69",
  1339 => x"74",
  1340 => x"0d",
  1341 => x"0a",
  1342 => x"00",
  1343 => x"49",
  1344 => x"6e",
  1345 => x"69",
  1346 => x"74",
  1347 => x"20",
  1348 => x"64",
  1349 => x"6f",
  1350 => x"6e",
  1351 => x"65",
  1352 => x"0d",
  1353 => x"0a",
  1354 => x"00",
  1355 => x"49",
  1356 => x"6e",
  1357 => x"69",
  1358 => x"74",
  1359 => x"20",
  1360 => x"66",
  1361 => x"61",
  1362 => x"69",
  1363 => x"6c",
  1364 => x"75",
  1365 => x"72",
  1366 => x"65",
  1367 => x"0d",
  1368 => x"0a",
  1369 => x"00",
  1370 => x"52",
  1371 => x"65",
  1372 => x"73",
  1373 => x"65",
  1374 => x"74",
  1375 => x"20",
  1376 => x"66",
  1377 => x"61",
  1378 => x"69",
  1379 => x"6c",
  1380 => x"75",
  1381 => x"72",
  1382 => x"65",
  1383 => x"0d",
  1384 => x"0a",
  1385 => x"00",
  1386 => x"43",
  1387 => x"6f",
  1388 => x"6d",
  1389 => x"6d",
  1390 => x"61",
  1391 => x"6e",
  1392 => x"64",
  1393 => x"20",
  1394 => x"54",
  1395 => x"69",
  1396 => x"6d",
  1397 => x"65",
  1398 => x"6f",
  1399 => x"75",
  1400 => x"74",
  1401 => x"5f",
  1402 => x"45",
  1403 => x"72",
  1404 => x"72",
  1405 => x"6f",
  1406 => x"72",
  1407 => x"0d",
  1408 => x"0a",
  1409 => x"00",
  1410 => x"54",
  1411 => x"69",
  1412 => x"6d",
  1413 => x"65",
  1414 => x"6f",
  1415 => x"75",
  1416 => x"74",
  1417 => x"5f",
  1418 => x"45",
  1419 => x"72",
  1420 => x"72",
  1421 => x"6f",
  1422 => x"72",
  1423 => x"0d",
  1424 => x"0a",
  1425 => x"00",
  1426 => x"53",
  1427 => x"44",
  1428 => x"48",
  1429 => x"43",
  1430 => x"20",
  1431 => x"66",
  1432 => x"6f",
  1433 => x"75",
  1434 => x"6e",
  1435 => x"64",
  1436 => x"20",
  1437 => x"0d",
  1438 => x"0a",
  1439 => x"00",
  1440 => x"33",
  1441 => x"fc",
  1442 => x"ff",
  1443 => x"ff",
  1444 => x"00",
  1445 => x"7f",
  1446 => x"00",
  1447 => x"24",
  1448 => x"43",
  1449 => x"f9",
  1450 => x"81",
  1451 => x"00",
  1452 => x"00",
  1453 => x"00",
  1454 => x"33",
  1455 => x"7c",
  1456 => x"00",
  1457 => x"00",
  1458 => x"00",
  1459 => x"22",
  1460 => x"33",
  1461 => x"7c",
  1462 => x"00",
  1463 => x"96",
  1464 => x"00",
  1465 => x"1e",
  1466 => x"32",
  1467 => x"3c",
  1468 => x"00",
  1469 => x"c8",
  1470 => x"43",
  1471 => x"e9",
  1472 => x"00",
  1473 => x"20",
  1474 => x"33",
  1475 => x"7c",
  1476 => x"00",
  1477 => x"ff",
  1478 => x"00",
  1479 => x"24",
  1480 => x"51",
  1481 => x"c9",
  1482 => x"ff",
  1483 => x"f8",
  1484 => x"34",
  1485 => x"3c",
  1486 => x"00",
  1487 => x"32",
  1488 => x"61",
  1489 => x"00",
  1490 => x"fe",
  1491 => x"96",
  1492 => x"3f",
  1493 => x"69",
  1494 => x"00",
  1495 => x"24",
  1496 => x"ff",
  1497 => x"fe",
  1498 => x"33",
  1499 => x"7c",
  1500 => x"00",
  1501 => x"00",
  1502 => x"00",
  1503 => x"22",
  1504 => x"b0",
  1505 => x"3c",
  1506 => x"00",
  1507 => x"01",
  1508 => x"67",
  1509 => x"12",
  1510 => x"51",
  1511 => x"ca",
  1512 => x"ff",
  1513 => x"e8",
  1514 => x"48",
  1515 => x"7a",
  1516 => x"ff",
  1517 => x"6e",
  1518 => x"61",
  1519 => x"00",
  1520 => x"01",
  1521 => x"22",
  1522 => x"58",
  1523 => x"8f",
  1524 => x"70",
  1525 => x"ff",
  1526 => x"4e",
  1527 => x"75",
  1528 => x"22",
  1529 => x"3c",
  1530 => x"00",
  1531 => x"00",
  1532 => x"20",
  1533 => x"00",
  1534 => x"33",
  1535 => x"7c",
  1536 => x"00",
  1537 => x"ff",
  1538 => x"00",
  1539 => x"24",
  1540 => x"53",
  1541 => x"81",
  1542 => x"66",
  1543 => x"f6",
  1544 => x"61",
  1545 => x"00",
  1546 => x"fe",
  1547 => x"72",
  1548 => x"b0",
  1549 => x"3c",
  1550 => x"00",
  1551 => x"01",
  1552 => x"66",
  1553 => x"00",
  1554 => x"00",
  1555 => x"9e",
  1556 => x"33",
  1557 => x"7c",
  1558 => x"00",
  1559 => x"ff",
  1560 => x"00",
  1561 => x"24",
  1562 => x"33",
  1563 => x"7c",
  1564 => x"00",
  1565 => x"ff",
  1566 => x"00",
  1567 => x"24",
  1568 => x"33",
  1569 => x"7c",
  1570 => x"00",
  1571 => x"ff",
  1572 => x"00",
  1573 => x"24",
  1574 => x"30",
  1575 => x"29",
  1576 => x"00",
  1577 => x"24",
  1578 => x"0c",
  1579 => x"00",
  1580 => x"00",
  1581 => x"01",
  1582 => x"66",
  1583 => x"00",
  1584 => x"00",
  1585 => x"80",
  1586 => x"33",
  1587 => x"7c",
  1588 => x"00",
  1589 => x"ff",
  1590 => x"00",
  1591 => x"24",
  1592 => x"30",
  1593 => x"29",
  1594 => x"00",
  1595 => x"24",
  1596 => x"0c",
  1597 => x"00",
  1598 => x"00",
  1599 => x"aa",
  1600 => x"66",
  1601 => x"6e",
  1602 => x"3f",
  1603 => x"69",
  1604 => x"00",
  1605 => x"24",
  1606 => x"ff",
  1607 => x"fe",
  1608 => x"33",
  1609 => x"7c",
  1610 => x"00",
  1611 => x"00",
  1612 => x"00",
  1613 => x"22",
  1614 => x"48",
  1615 => x"7a",
  1616 => x"ff",
  1617 => x"42",
  1618 => x"61",
  1619 => x"00",
  1620 => x"00",
  1621 => x"be",
  1622 => x"58",
  1623 => x"8f",
  1624 => x"34",
  1625 => x"3c",
  1626 => x"00",
  1627 => x"32",
  1628 => x"53",
  1629 => x"42",
  1630 => x"67",
  1631 => x"50",
  1632 => x"32",
  1633 => x"3c",
  1634 => x"07",
  1635 => x"d0",
  1636 => x"33",
  1637 => x"7c",
  1638 => x"00",
  1639 => x"ff",
  1640 => x"00",
  1641 => x"24",
  1642 => x"51",
  1643 => x"c9",
  1644 => x"ff",
  1645 => x"f8",
  1646 => x"61",
  1647 => x"00",
  1648 => x"fe",
  1649 => x"28",
  1650 => x"b0",
  1651 => x"3c",
  1652 => x"00",
  1653 => x"01",
  1654 => x"66",
  1655 => x"e4",
  1656 => x"61",
  1657 => x"00",
  1658 => x"fe",
  1659 => x"10",
  1660 => x"66",
  1661 => x"de",
  1662 => x"61",
  1663 => x"00",
  1664 => x"fe",
  1665 => x"22",
  1666 => x"66",
  1667 => x"d8",
  1668 => x"33",
  1669 => x"7c",
  1670 => x"00",
  1671 => x"ff",
  1672 => x"00",
  1673 => x"24",
  1674 => x"30",
  1675 => x"29",
  1676 => x"00",
  1677 => x"24",
  1678 => x"c0",
  1679 => x"3c",
  1680 => x"00",
  1681 => x"40",
  1682 => x"66",
  1683 => x"08",
  1684 => x"33",
  1685 => x"fc",
  1686 => x"00",
  1687 => x"00",
  1688 => x"00",
  1689 => x"7f",
  1690 => x"00",
  1691 => x"24",
  1692 => x"33",
  1693 => x"7c",
  1694 => x"00",
  1695 => x"ff",
  1696 => x"00",
  1697 => x"24",
  1698 => x"33",
  1699 => x"7c",
  1700 => x"00",
  1701 => x"ff",
  1702 => x"00",
  1703 => x"24",
  1704 => x"33",
  1705 => x"7c",
  1706 => x"00",
  1707 => x"ff",
  1708 => x"00",
  1709 => x"24",
  1710 => x"60",
  1711 => x"3c",
  1712 => x"33",
  1713 => x"fc",
  1714 => x"00",
  1715 => x"00",
  1716 => x"00",
  1717 => x"7f",
  1718 => x"00",
  1719 => x"24",
  1720 => x"34",
  1721 => x"3c",
  1722 => x"00",
  1723 => x"0a",
  1724 => x"32",
  1725 => x"3c",
  1726 => x"07",
  1727 => x"d0",
  1728 => x"33",
  1729 => x"7c",
  1730 => x"00",
  1731 => x"ff",
  1732 => x"00",
  1733 => x"24",
  1734 => x"51",
  1735 => x"c9",
  1736 => x"ff",
  1737 => x"f8",
  1738 => x"61",
  1739 => x"00",
  1740 => x"fd",
  1741 => x"a6",
  1742 => x"67",
  1743 => x"1c",
  1744 => x"3f",
  1745 => x"69",
  1746 => x"00",
  1747 => x"24",
  1748 => x"ff",
  1749 => x"fe",
  1750 => x"33",
  1751 => x"7c",
  1752 => x"00",
  1753 => x"00",
  1754 => x"00",
  1755 => x"22",
  1756 => x"51",
  1757 => x"ca",
  1758 => x"ff",
  1759 => x"de",
  1760 => x"48",
  1761 => x"7a",
  1762 => x"fe",
  1763 => x"69",
  1764 => x"61",
  1765 => x"2c",
  1766 => x"58",
  1767 => x"8f",
  1768 => x"70",
  1769 => x"ff",
  1770 => x"4e",
  1771 => x"75",
  1772 => x"3f",
  1773 => x"69",
  1774 => x"00",
  1775 => x"24",
  1776 => x"ff",
  1777 => x"fe",
  1778 => x"33",
  1779 => x"7c",
  1780 => x"00",
  1781 => x"00",
  1782 => x"00",
  1783 => x"22",
  1784 => x"33",
  1785 => x"69",
  1786 => x"00",
  1787 => x"2c",
  1788 => x"00",
  1789 => x"1e",
  1790 => x"48",
  1791 => x"7a",
  1792 => x"fe",
  1793 => x"3f",
  1794 => x"61",
  1795 => x"0e",
  1796 => x"58",
  1797 => x"8f",
  1798 => x"33",
  1799 => x"fc",
  1800 => x"ff",
  1801 => x"ff",
  1802 => x"81",
  1803 => x"00",
  1804 => x"00",
  1805 => x"06",
  1806 => x"70",
  1807 => x"00",
  1808 => x"4e",
  1809 => x"75",
  1810 => x"2f",
  1811 => x"08",
  1812 => x"20",
  1813 => x"6f",
  1814 => x"00",
  1815 => x"08",
  1816 => x"61",
  1817 => x"04",
  1818 => x"20",
  1819 => x"5f",
  1820 => x"4e",
  1821 => x"75",
  1822 => x"48",
  1823 => x"e7",
  1824 => x"00",
  1825 => x"c0",
  1826 => x"22",
  1827 => x"39",
  1828 => x"00",
  1829 => x"7f",
  1830 => x"00",
  1831 => x"52",
  1832 => x"43",
  1833 => x"f9",
  1834 => x"80",
  1835 => x"00",
  1836 => x"08",
  1837 => x"00",
  1838 => x"10",
  1839 => x"18",
  1840 => x"67",
  1841 => x"08",
  1842 => x"13",
  1843 => x"80",
  1844 => x"10",
  1845 => x"00",
  1846 => x"52",
  1847 => x"41",
  1848 => x"60",
  1849 => x"f4",
  1850 => x"06",
  1851 => x"b9",
  1852 => x"00",
  1853 => x"00",
  1854 => x"00",
  1855 => x"4c",
  1856 => x"00",
  1857 => x"7f",
  1858 => x"00",
  1859 => x"52",
  1860 => x"4c",
  1861 => x"df",
  1862 => x"03",
  1863 => x"00",
  1864 => x"4e",
  1865 => x"75",
  1866 => x"4a",
  1867 => x"79",
  1868 => x"00",
  1869 => x"7f",
  1870 => x"00",
  1871 => x"24",
  1872 => x"67",
  1873 => x"1e",
  1874 => x"41",
  1875 => x"fa",
  1876 => x"00",
  1877 => x"08",
  1878 => x"48",
  1879 => x"7a",
  1880 => x"00",
  1881 => x"34",
  1882 => x"60",
  1883 => x"c2",
  1884 => x"53",
  1885 => x"44",
  1886 => x"48",
  1887 => x"43",
  1888 => x"20",
  1889 => x"66",
  1890 => x"6c",
  1891 => x"61",
  1892 => x"67",
  1893 => x"20",
  1894 => x"73",
  1895 => x"74",
  1896 => x"69",
  1897 => x"6c",
  1898 => x"6c",
  1899 => x"20",
  1900 => x"73",
  1901 => x"65",
  1902 => x"74",
  1903 => x"00",
  1904 => x"41",
  1905 => x"fa",
  1906 => x"00",
  1907 => x"08",
  1908 => x"48",
  1909 => x"7a",
  1910 => x"00",
  1911 => x"16",
  1912 => x"60",
  1913 => x"a4",
  1914 => x"53",
  1915 => x"44",
  1916 => x"48",
  1917 => x"43",
  1918 => x"20",
  1919 => x"66",
  1920 => x"6c",
  1921 => x"61",
  1922 => x"67",
  1923 => x"20",
  1924 => x"63",
  1925 => x"6c",
  1926 => x"65",
  1927 => x"61",
  1928 => x"72",
  1929 => x"65",
  1930 => x"64",
  1931 => x"00",
  1932 => x"61",
  1933 => x"00",
  1934 => x"02",
  1935 => x"0a",
  1936 => x"61",
  1937 => x"00",
  1938 => x"fc",
  1939 => x"46",
  1940 => x"66",
  1941 => x"46",
  1942 => x"2e",
  1943 => x"3c",
  1944 => x"00",
  1945 => x"00",
  1946 => x"01",
  1947 => x"ff",
  1948 => x"41",
  1949 => x"f9",
  1950 => x"00",
  1951 => x"7f",
  1952 => x"00",
  1953 => x"56",
  1954 => x"43",
  1955 => x"f9",
  1956 => x"80",
  1957 => x"00",
  1958 => x"08",
  1959 => x"00",
  1960 => x"10",
  1961 => x"18",
  1962 => x"12",
  1963 => x"c0",
  1964 => x"48",
  1965 => x"e7",
  1966 => x"01",
  1967 => x"c0",
  1968 => x"61",
  1969 => x"00",
  1970 => x"f9",
  1971 => x"70",
  1972 => x"4c",
  1973 => x"df",
  1974 => x"03",
  1975 => x"80",
  1976 => x"51",
  1977 => x"cf",
  1978 => x"ff",
  1979 => x"ee",
  1980 => x"20",
  1981 => x"39",
  1982 => x"00",
  1983 => x"7f",
  1984 => x"00",
  1985 => x"38",
  1986 => x"52",
  1987 => x"80",
  1988 => x"23",
  1989 => x"c0",
  1990 => x"00",
  1991 => x"7f",
  1992 => x"00",
  1993 => x"38",
  1994 => x"53",
  1995 => x"79",
  1996 => x"00",
  1997 => x"7f",
  1998 => x"00",
  1999 => x"36",
  2000 => x"66",
  2001 => x"be",
  2002 => x"61",
  2003 => x"00",
  2004 => x"02",
  2005 => x"7a",
  2006 => x"66",
  2007 => x"b4",
  2008 => x"20",
  2009 => x"08",
  2010 => x"4e",
  2011 => x"75",
  2012 => x"70",
  2013 => x"00",
  2014 => x"4e",
  2015 => x"75",
  2016 => x"33",
  2017 => x"fc",
  2018 => x"02",
  2019 => x"01",
  2020 => x"81",
  2021 => x"00",
  2022 => x"00",
  2023 => x"06",
  2024 => x"70",
  2025 => x"00",
  2026 => x"23",
  2027 => x"c0",
  2028 => x"00",
  2029 => x"7f",
  2030 => x"00",
  2031 => x"3e",
  2032 => x"33",
  2033 => x"fc",
  2034 => x"02",
  2035 => x"11",
  2036 => x"81",
  2037 => x"00",
  2038 => x"00",
  2039 => x"06",
  2040 => x"61",
  2041 => x"00",
  2042 => x"fb",
  2043 => x"de",
  2044 => x"66",
  2045 => x"5c",
  2046 => x"33",
  2047 => x"fc",
  2048 => x"02",
  2049 => x"02",
  2050 => x"81",
  2051 => x"00",
  2052 => x"00",
  2053 => x"06",
  2054 => x"0c",
  2055 => x"28",
  2056 => x"00",
  2057 => x"55",
  2058 => x"01",
  2059 => x"fe",
  2060 => x"66",
  2061 => x"4c",
  2062 => x"0c",
  2063 => x"28",
  2064 => x"00",
  2065 => x"aa",
  2066 => x"01",
  2067 => x"ff",
  2068 => x"66",
  2069 => x"44",
  2070 => x"30",
  2071 => x"39",
  2072 => x"00",
  2073 => x"7f",
  2074 => x"00",
  2075 => x"26",
  2076 => x"c0",
  2077 => x"7c",
  2078 => x"00",
  2079 => x"70",
  2080 => x"b0",
  2081 => x"7c",
  2082 => x"00",
  2083 => x"40",
  2084 => x"64",
  2085 => x"40",
  2086 => x"43",
  2087 => x"e8",
  2088 => x"01",
  2089 => x"be",
  2090 => x"d2",
  2091 => x"c0",
  2092 => x"33",
  2093 => x"fc",
  2094 => x"02",
  2095 => x"03",
  2096 => x"81",
  2097 => x"00",
  2098 => x"00",
  2099 => x"06",
  2100 => x"20",
  2101 => x"29",
  2102 => x"00",
  2103 => x"08",
  2104 => x"e0",
  2105 => x"58",
  2106 => x"48",
  2107 => x"40",
  2108 => x"e0",
  2109 => x"58",
  2110 => x"23",
  2111 => x"c0",
  2112 => x"00",
  2113 => x"7f",
  2114 => x"00",
  2115 => x"3e",
  2116 => x"61",
  2117 => x"00",
  2118 => x"fb",
  2119 => x"92",
  2120 => x"66",
  2121 => x"10",
  2122 => x"0c",
  2123 => x"28",
  2124 => x"00",
  2125 => x"55",
  2126 => x"01",
  2127 => x"fe",
  2128 => x"66",
  2129 => x"08",
  2130 => x"0c",
  2131 => x"28",
  2132 => x"00",
  2133 => x"aa",
  2134 => x"01",
  2135 => x"ff",
  2136 => x"67",
  2137 => x"0c",
  2138 => x"33",
  2139 => x"fc",
  2140 => x"f2",
  2141 => x"01",
  2142 => x"81",
  2143 => x"00",
  2144 => x"00",
  2145 => x"06",
  2146 => x"70",
  2147 => x"ff",
  2148 => x"4e",
  2149 => x"75",
  2150 => x"33",
  2151 => x"fc",
  2152 => x"02",
  2153 => x"04",
  2154 => x"81",
  2155 => x"00",
  2156 => x"00",
  2157 => x"06",
  2158 => x"0c",
  2159 => x"a8",
  2160 => x"46",
  2161 => x"41",
  2162 => x"54",
  2163 => x"31",
  2164 => x"00",
  2165 => x"36",
  2166 => x"66",
  2167 => x"24",
  2168 => x"13",
  2169 => x"fc",
  2170 => x"00",
  2171 => x"0c",
  2172 => x"00",
  2173 => x"7f",
  2174 => x"00",
  2175 => x"28",
  2176 => x"0c",
  2177 => x"a8",
  2178 => x"32",
  2179 => x"20",
  2180 => x"20",
  2181 => x"20",
  2182 => x"00",
  2183 => x"3a",
  2184 => x"67",
  2185 => x"36",
  2186 => x"13",
  2187 => x"fc",
  2188 => x"00",
  2189 => x"10",
  2190 => x"00",
  2191 => x"7f",
  2192 => x"00",
  2193 => x"28",
  2194 => x"0c",
  2195 => x"a8",
  2196 => x"36",
  2197 => x"20",
  2198 => x"20",
  2199 => x"20",
  2200 => x"00",
  2201 => x"3a",
  2202 => x"67",
  2203 => x"24",
  2204 => x"13",
  2205 => x"fc",
  2206 => x"00",
  2207 => x"00",
  2208 => x"00",
  2209 => x"7f",
  2210 => x"00",
  2211 => x"28",
  2212 => x"0c",
  2213 => x"a8",
  2214 => x"46",
  2215 => x"41",
  2216 => x"54",
  2217 => x"33",
  2218 => x"00",
  2219 => x"52",
  2220 => x"66",
  2221 => x"ac",
  2222 => x"0c",
  2223 => x"a8",
  2224 => x"32",
  2225 => x"20",
  2226 => x"20",
  2227 => x"20",
  2228 => x"00",
  2229 => x"56",
  2230 => x"66",
  2231 => x"a2",
  2232 => x"13",
  2233 => x"fc",
  2234 => x"00",
  2235 => x"20",
  2236 => x"00",
  2237 => x"7f",
  2238 => x"00",
  2239 => x"28",
  2240 => x"20",
  2241 => x"28",
  2242 => x"00",
  2243 => x"0a",
  2244 => x"c0",
  2245 => x"bc",
  2246 => x"00",
  2247 => x"ff",
  2248 => x"ff",
  2249 => x"00",
  2250 => x"0c",
  2251 => x"80",
  2252 => x"00",
  2253 => x"00",
  2254 => x"02",
  2255 => x"00",
  2256 => x"66",
  2257 => x"88",
  2258 => x"22",
  2259 => x"39",
  2260 => x"00",
  2261 => x"7f",
  2262 => x"00",
  2263 => x"3e",
  2264 => x"30",
  2265 => x"28",
  2266 => x"00",
  2267 => x"0e",
  2268 => x"e0",
  2269 => x"58",
  2270 => x"d2",
  2271 => x"80",
  2272 => x"23",
  2273 => x"c1",
  2274 => x"00",
  2275 => x"7f",
  2276 => x"00",
  2277 => x"42",
  2278 => x"0c",
  2279 => x"39",
  2280 => x"00",
  2281 => x"20",
  2282 => x"00",
  2283 => x"7f",
  2284 => x"00",
  2285 => x"28",
  2286 => x"66",
  2287 => x"24",
  2288 => x"20",
  2289 => x"28",
  2290 => x"00",
  2291 => x"2c",
  2292 => x"e0",
  2293 => x"58",
  2294 => x"48",
  2295 => x"40",
  2296 => x"e0",
  2297 => x"58",
  2298 => x"23",
  2299 => x"c0",
  2300 => x"00",
  2301 => x"7f",
  2302 => x"00",
  2303 => x"2a",
  2304 => x"20",
  2305 => x"28",
  2306 => x"00",
  2307 => x"24",
  2308 => x"e0",
  2309 => x"58",
  2310 => x"48",
  2311 => x"40",
  2312 => x"e0",
  2313 => x"58",
  2314 => x"d2",
  2315 => x"80",
  2316 => x"53",
  2317 => x"28",
  2318 => x"00",
  2319 => x"10",
  2320 => x"66",
  2321 => x"f8",
  2322 => x"60",
  2323 => x"32",
  2324 => x"70",
  2325 => x"00",
  2326 => x"23",
  2327 => x"c0",
  2328 => x"00",
  2329 => x"7f",
  2330 => x"00",
  2331 => x"2a",
  2332 => x"30",
  2333 => x"28",
  2334 => x"00",
  2335 => x"16",
  2336 => x"e0",
  2337 => x"58",
  2338 => x"d2",
  2339 => x"80",
  2340 => x"53",
  2341 => x"28",
  2342 => x"00",
  2343 => x"10",
  2344 => x"66",
  2345 => x"f8",
  2346 => x"23",
  2347 => x"c1",
  2348 => x"00",
  2349 => x"7f",
  2350 => x"00",
  2351 => x"2e",
  2352 => x"20",
  2353 => x"01",
  2354 => x"10",
  2355 => x"28",
  2356 => x"00",
  2357 => x"12",
  2358 => x"e1",
  2359 => x"48",
  2360 => x"10",
  2361 => x"28",
  2362 => x"00",
  2363 => x"11",
  2364 => x"33",
  2365 => x"c0",
  2366 => x"00",
  2367 => x"7f",
  2368 => x"00",
  2369 => x"4e",
  2370 => x"e8",
  2371 => x"48",
  2372 => x"d2",
  2373 => x"80",
  2374 => x"70",
  2375 => x"00",
  2376 => x"10",
  2377 => x"28",
  2378 => x"00",
  2379 => x"0d",
  2380 => x"33",
  2381 => x"c0",
  2382 => x"00",
  2383 => x"7f",
  2384 => x"00",
  2385 => x"4a",
  2386 => x"92",
  2387 => x"80",
  2388 => x"92",
  2389 => x"80",
  2390 => x"23",
  2391 => x"c1",
  2392 => x"00",
  2393 => x"7f",
  2394 => x"00",
  2395 => x"46",
  2396 => x"33",
  2397 => x"fc",
  2398 => x"02",
  2399 => x"05",
  2400 => x"81",
  2401 => x"00",
  2402 => x"00",
  2403 => x"06",
  2404 => x"70",
  2405 => x"00",
  2406 => x"4e",
  2407 => x"75",
  2408 => x"20",
  2409 => x"39",
  2410 => x"00",
  2411 => x"7f",
  2412 => x"00",
  2413 => x"2a",
  2414 => x"23",
  2415 => x"c0",
  2416 => x"00",
  2417 => x"7f",
  2418 => x"00",
  2419 => x"32",
  2420 => x"66",
  2421 => x"28",
  2422 => x"42",
  2423 => x"b9",
  2424 => x"00",
  2425 => x"7f",
  2426 => x"00",
  2427 => x"32",
  2428 => x"30",
  2429 => x"39",
  2430 => x"00",
  2431 => x"7f",
  2432 => x"00",
  2433 => x"4e",
  2434 => x"e8",
  2435 => x"48",
  2436 => x"33",
  2437 => x"c0",
  2438 => x"00",
  2439 => x"7f",
  2440 => x"00",
  2441 => x"36",
  2442 => x"20",
  2443 => x"39",
  2444 => x"00",
  2445 => x"7f",
  2446 => x"00",
  2447 => x"2e",
  2448 => x"23",
  2449 => x"c0",
  2450 => x"00",
  2451 => x"7f",
  2452 => x"00",
  2453 => x"38",
  2454 => x"4e",
  2455 => x"75",
  2456 => x"20",
  2457 => x"39",
  2458 => x"00",
  2459 => x"7f",
  2460 => x"00",
  2461 => x"32",
  2462 => x"32",
  2463 => x"39",
  2464 => x"00",
  2465 => x"7f",
  2466 => x"00",
  2467 => x"4a",
  2468 => x"33",
  2469 => x"c1",
  2470 => x"00",
  2471 => x"7f",
  2472 => x"00",
  2473 => x"36",
  2474 => x"e2",
  2475 => x"49",
  2476 => x"65",
  2477 => x"04",
  2478 => x"e3",
  2479 => x"88",
  2480 => x"60",
  2481 => x"f8",
  2482 => x"d0",
  2483 => x"b9",
  2484 => x"00",
  2485 => x"7f",
  2486 => x"00",
  2487 => x"46",
  2488 => x"23",
  2489 => x"c0",
  2490 => x"00",
  2491 => x"7f",
  2492 => x"00",
  2493 => x"38",
  2494 => x"4e",
  2495 => x"75",
  2496 => x"48",
  2497 => x"e7",
  2498 => x"20",
  2499 => x"20",
  2500 => x"24",
  2501 => x"49",
  2502 => x"61",
  2503 => x"00",
  2504 => x"fa",
  2505 => x"10",
  2506 => x"66",
  2507 => x"7a",
  2508 => x"74",
  2509 => x"0f",
  2510 => x"4a",
  2511 => x"10",
  2512 => x"67",
  2513 => x"74",
  2514 => x"70",
  2515 => x"0a",
  2516 => x"12",
  2517 => x"32",
  2518 => x"00",
  2519 => x"00",
  2520 => x"b2",
  2521 => x"30",
  2522 => x"00",
  2523 => x"00",
  2524 => x"67",
  2525 => x"0a",
  2526 => x"d2",
  2527 => x"3c",
  2528 => x"00",
  2529 => x"20",
  2530 => x"b2",
  2531 => x"30",
  2532 => x"00",
  2533 => x"00",
  2534 => x"66",
  2535 => x"36",
  2536 => x"51",
  2537 => x"c8",
  2538 => x"ff",
  2539 => x"ea",
  2540 => x"70",
  2541 => x"00",
  2542 => x"10",
  2543 => x"28",
  2544 => x"00",
  2545 => x"0b",
  2546 => x"33",
  2547 => x"c0",
  2548 => x"00",
  2549 => x"7f",
  2550 => x"00",
  2551 => x"3c",
  2552 => x"0c",
  2553 => x"39",
  2554 => x"00",
  2555 => x"20",
  2556 => x"00",
  2557 => x"7f",
  2558 => x"00",
  2559 => x"28",
  2560 => x"66",
  2561 => x"08",
  2562 => x"30",
  2563 => x"28",
  2564 => x"00",
  2565 => x"14",
  2566 => x"e0",
  2567 => x"58",
  2568 => x"48",
  2569 => x"40",
  2570 => x"30",
  2571 => x"28",
  2572 => x"00",
  2573 => x"1a",
  2574 => x"e0",
  2575 => x"58",
  2576 => x"23",
  2577 => x"c0",
  2578 => x"00",
  2579 => x"7f",
  2580 => x"00",
  2581 => x"32",
  2582 => x"4c",
  2583 => x"df",
  2584 => x"04",
  2585 => x"04",
  2586 => x"70",
  2587 => x"ff",
  2588 => x"4e",
  2589 => x"75",
  2590 => x"41",
  2591 => x"e8",
  2592 => x"00",
  2593 => x"20",
  2594 => x"51",
  2595 => x"ca",
  2596 => x"ff",
  2597 => x"aa",
  2598 => x"20",
  2599 => x"39",
  2600 => x"00",
  2601 => x"7f",
  2602 => x"00",
  2603 => x"38",
  2604 => x"52",
  2605 => x"80",
  2606 => x"23",
  2607 => x"c0",
  2608 => x"00",
  2609 => x"7f",
  2610 => x"00",
  2611 => x"38",
  2612 => x"53",
  2613 => x"79",
  2614 => x"00",
  2615 => x"7f",
  2616 => x"00",
  2617 => x"36",
  2618 => x"66",
  2619 => x"8a",
  2620 => x"61",
  2621 => x"10",
  2622 => x"67",
  2623 => x"06",
  2624 => x"61",
  2625 => x"00",
  2626 => x"ff",
  2627 => x"56",
  2628 => x"60",
  2629 => x"80",
  2630 => x"4c",
  2631 => x"df",
  2632 => x"04",
  2633 => x"04",
  2634 => x"70",
  2635 => x"00",
  2636 => x"4e",
  2637 => x"75",
  2638 => x"0c",
  2639 => x"39",
  2640 => x"00",
  2641 => x"20",
  2642 => x"00",
  2643 => x"7f",
  2644 => x"00",
  2645 => x"28",
  2646 => x"67",
  2647 => x"3e",
  2648 => x"0c",
  2649 => x"39",
  2650 => x"00",
  2651 => x"0c",
  2652 => x"00",
  2653 => x"7f",
  2654 => x"00",
  2655 => x"28",
  2656 => x"67",
  2657 => x"78",
  2658 => x"20",
  2659 => x"39",
  2660 => x"00",
  2661 => x"7f",
  2662 => x"00",
  2663 => x"32",
  2664 => x"e0",
  2665 => x"88",
  2666 => x"d0",
  2667 => x"b9",
  2668 => x"00",
  2669 => x"7f",
  2670 => x"00",
  2671 => x"42",
  2672 => x"61",
  2673 => x"00",
  2674 => x"f9",
  2675 => x"66",
  2676 => x"66",
  2677 => x"60",
  2678 => x"10",
  2679 => x"39",
  2680 => x"00",
  2681 => x"7f",
  2682 => x"00",
  2683 => x"35",
  2684 => x"d0",
  2685 => x"40",
  2686 => x"30",
  2687 => x"30",
  2688 => x"00",
  2689 => x"00",
  2690 => x"e0",
  2691 => x"58",
  2692 => x"23",
  2693 => x"c0",
  2694 => x"00",
  2695 => x"7f",
  2696 => x"00",
  2697 => x"32",
  2698 => x"80",
  2699 => x"bc",
  2700 => x"ff",
  2701 => x"ff",
  2702 => x"00",
  2703 => x"0f",
  2704 => x"b0",
  2705 => x"7c",
  2706 => x"ff",
  2707 => x"ff",
  2708 => x"4e",
  2709 => x"75",
  2710 => x"20",
  2711 => x"39",
  2712 => x"00",
  2713 => x"7f",
  2714 => x"00",
  2715 => x"32",
  2716 => x"ee",
  2717 => x"88",
  2718 => x"d0",
  2719 => x"b9",
  2720 => x"00",
  2721 => x"7f",
  2722 => x"00",
  2723 => x"42",
  2724 => x"61",
  2725 => x"00",
  2726 => x"f9",
  2727 => x"32",
  2728 => x"66",
  2729 => x"2c",
  2730 => x"10",
  2731 => x"39",
  2732 => x"00",
  2733 => x"7f",
  2734 => x"00",
  2735 => x"35",
  2736 => x"c0",
  2737 => x"7c",
  2738 => x"00",
  2739 => x"7f",
  2740 => x"d0",
  2741 => x"40",
  2742 => x"d0",
  2743 => x"40",
  2744 => x"20",
  2745 => x"30",
  2746 => x"00",
  2747 => x"00",
  2748 => x"e0",
  2749 => x"58",
  2750 => x"48",
  2751 => x"40",
  2752 => x"e0",
  2753 => x"58",
  2754 => x"23",
  2755 => x"c0",
  2756 => x"00",
  2757 => x"7f",
  2758 => x"00",
  2759 => x"32",
  2760 => x"80",
  2761 => x"bc",
  2762 => x"f0",
  2763 => x"00",
  2764 => x"00",
  2765 => x"07",
  2766 => x"b0",
  2767 => x"bc",
  2768 => x"ff",
  2769 => x"ff",
  2770 => x"ff",
  2771 => x"ff",
  2772 => x"4e",
  2773 => x"75",
  2774 => x"70",
  2775 => x"00",
  2776 => x"4e",
  2777 => x"75",
  2778 => x"2f",
  2779 => x"02",
  2780 => x"20",
  2781 => x"39",
  2782 => x"00",
  2783 => x"7f",
  2784 => x"00",
  2785 => x"32",
  2786 => x"22",
  2787 => x"00",
  2788 => x"d0",
  2789 => x"80",
  2790 => x"d0",
  2791 => x"81",
  2792 => x"22",
  2793 => x"00",
  2794 => x"e0",
  2795 => x"88",
  2796 => x"e4",
  2797 => x"88",
  2798 => x"d0",
  2799 => x"b9",
  2800 => x"00",
  2801 => x"7f",
  2802 => x"00",
  2803 => x"42",
  2804 => x"24",
  2805 => x"00",
  2806 => x"61",
  2807 => x"00",
  2808 => x"f8",
  2809 => x"e0",
  2810 => x"66",
  2811 => x"52",
  2812 => x"20",
  2813 => x"01",
  2814 => x"e2",
  2815 => x"88",
  2816 => x"c0",
  2817 => x"7c",
  2818 => x"01",
  2819 => x"ff",
  2820 => x"b0",
  2821 => x"7c",
  2822 => x"01",
  2823 => x"ff",
  2824 => x"66",
  2825 => x"14",
  2826 => x"10",
  2827 => x"30",
  2828 => x"00",
  2829 => x"00",
  2830 => x"c1",
  2831 => x"42",
  2832 => x"52",
  2833 => x"80",
  2834 => x"61",
  2835 => x"00",
  2836 => x"f8",
  2837 => x"c4",
  2838 => x"66",
  2839 => x"36",
  2840 => x"e1",
  2841 => x"4a",
  2842 => x"14",
  2843 => x"10",
  2844 => x"60",
  2845 => x"0a",
  2846 => x"14",
  2847 => x"30",
  2848 => x"00",
  2849 => x"00",
  2850 => x"e1",
  2851 => x"4a",
  2852 => x"14",
  2853 => x"30",
  2854 => x"00",
  2855 => x"01",
  2856 => x"e1",
  2857 => x"5a",
  2858 => x"c2",
  2859 => x"7c",
  2860 => x"00",
  2861 => x"01",
  2862 => x"67",
  2863 => x"02",
  2864 => x"e8",
  2865 => x"4a",
  2866 => x"c4",
  2867 => x"bc",
  2868 => x"00",
  2869 => x"00",
  2870 => x"0f",
  2871 => x"ff",
  2872 => x"23",
  2873 => x"c2",
  2874 => x"00",
  2875 => x"7f",
  2876 => x"00",
  2877 => x"32",
  2878 => x"84",
  2879 => x"bc",
  2880 => x"ff",
  2881 => x"ff",
  2882 => x"f0",
  2883 => x"0f",
  2884 => x"20",
  2885 => x"02",
  2886 => x"24",
  2887 => x"1f",
  2888 => x"b0",
  2889 => x"7c",
  2890 => x"ff",
  2891 => x"ff",
  2892 => x"4e",
  2893 => x"75",
  2894 => x"24",
  2895 => x"1f",
  2896 => x"70",
  2897 => x"00",
  2898 => x"4e",
  2899 => x"75",
  2900 => x"41",
  2901 => x"f9",
  2902 => x"00",
  2903 => x"7f",
  2904 => x"00",
  2905 => x"04",
  2906 => x"20",
  2907 => x"bc",
  2908 => x"12",
  2909 => x"34",
  2910 => x"56",
  2911 => x"78",
  2912 => x"21",
  2913 => x"7c",
  2914 => x"fe",
  2915 => x"dc",
  2916 => x"ba",
  2917 => x"98",
  2918 => x"00",
  2919 => x"04",
  2920 => x"21",
  2921 => x"7c",
  2922 => x"aa",
  2923 => x"55",
  2924 => x"cc",
  2925 => x"22",
  2926 => x"00",
  2927 => x"02",
  2928 => x"11",
  2929 => x"7c",
  2930 => x"00",
  2931 => x"33",
  2932 => x"00",
  2933 => x"03",
  2934 => x"11",
  2935 => x"7c",
  2936 => x"00",
  2937 => x"fe",
  2938 => x"00",
  2939 => x"04",
  2940 => x"20",
  2941 => x"10",
  2942 => x"22",
  2943 => x"28",
  2944 => x"00",
  2945 => x"04",
  2946 => x"90",
  2947 => x"bc",
  2948 => x"12",
  2949 => x"34",
  2950 => x"aa",
  2951 => x"33",
  2952 => x"92",
  2953 => x"bc",
  2954 => x"fe",
  2955 => x"22",
  2956 => x"ba",
  2957 => x"98",
  2958 => x"80",
  2959 => x"81",
  2960 => x"4e",
  2961 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity video_vga_dither is
	port (
		pixelclock : in std_logic;
		X : in unsigned(9 downto 0);
		Y : in unsigned(9 downto 0);
		VSync : in std_logic;
		enable : in std_logic;
		iRed : in unsigned(7 downto 0);
		iGreen : in unsigned(7 downto 0);
		iBlue : in unsigned(7 downto 0);
		oRed : out unsigned(3 downto 0);
		oGreen : out unsigned(3 downto 0);
		oBlue : out unsigned(3 downto 0)
	);
end entity;

architecture rtl of video_vga_dither is
	signal field : std_logic := '0';
	signal red : unsigned(7 downto 0);
	signal green : unsigned(7 downto 0);
	signal blue : unsigned(7 downto 0);
begin

	oRed <= red(7 downto 4);
	oGreen <= green(7 downto 4);
	oBlue <= blue(7 downto 4);

	process(VSync,field)
	begin
		if rising_edge(VSync) then
			field <= not field;
		end if;
	end process;
	
	process(pixelclock,iRed,iGreen,iBlue,X,Y,field)
	begin
		if(rising_edge(pixelclock)) then
		
			if iRed(7 downto 4)="1111" or enable='0' then
				red <= iRed;
			else
				red <= (iRed + ((field xor Y(0)) & (X(0) xor Y(0)) & "00"));
			end if;
			
			if iGreen(7 downto 4)="1111" or enable='0' then
				green <= iGreen;
			else
				green <= (iGreen + ((field xor Y(0)) & (X(0) xor Y(0)) & "00"));
			end if;

			if iBlue(7 downto 4)="1111" or enable='0' then
				blue <= iBlue;
			else
				blue <= (iBlue+ ((field xor Y(0)) & (X(0) xor Y(0)) & "00"));
			end if;
			
		end if;
	end process;
end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"41",
    49 => x"fa",
    50 => x"00",
    51 => x"72",
    52 => x"61",
    53 => x"00",
    54 => x"02",
    55 => x"d6",
    56 => x"33",
    57 => x"fc",
    58 => x"0f",
    59 => x"00",
    60 => x"81",
    61 => x"00",
    62 => x"00",
    63 => x"06",
    64 => x"2e",
    65 => x"3c",
    66 => x"00",
    67 => x"00",
    68 => x"07",
    69 => x"ff",
    70 => x"41",
    71 => x"f9",
    72 => x"80",
    73 => x"00",
    74 => x"08",
    75 => x"00",
    76 => x"10",
    77 => x"fc",
    78 => x"00",
    79 => x"20",
    80 => x"51",
    81 => x"cf",
    82 => x"ff",
    83 => x"fa",
    84 => x"23",
    85 => x"fc",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"7f",
    92 => x"00",
    93 => x"52",
    94 => x"41",
    95 => x"fa",
    96 => x"00",
    97 => x"44",
    98 => x"61",
    99 => x"00",
   100 => x"06",
   101 => x"b8",
   102 => x"61",
   103 => x"00",
   104 => x"0a",
   105 => x"ea",
   106 => x"4a",
   107 => x"80",
   108 => x"67",
   109 => x"0a",
   110 => x"41",
   111 => x"fa",
   112 => x"00",
   113 => x"68",
   114 => x"61",
   115 => x"00",
   116 => x"06",
   117 => x"a8",
   118 => x"60",
   119 => x"fe",
   120 => x"41",
   121 => x"fa",
   122 => x"00",
   123 => x"47",
   124 => x"61",
   125 => x"00",
   126 => x"06",
   127 => x"9e",
   128 => x"61",
   129 => x"00",
   130 => x"02",
   131 => x"aa",
   132 => x"4b",
   133 => x"f9",
   134 => x"80",
   135 => x"00",
   136 => x"08",
   137 => x"00",
   138 => x"33",
   139 => x"fc",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"7f",
   144 => x"00",
   145 => x"0c",
   146 => x"30",
   147 => x"39",
   148 => x"81",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"08",
   153 => x"00",
   154 => x"00",
   155 => x"09",
   156 => x"67",
   157 => x"f4",
   158 => x"1a",
   159 => x"c0",
   160 => x"61",
   161 => x"7e",
   162 => x"60",
   163 => x"ee",
   164 => x"43",
   165 => x"6f",
   166 => x"6e",
   167 => x"64",
   168 => x"75",
   169 => x"63",
   170 => x"74",
   171 => x"69",
   172 => x"6e",
   173 => x"67",
   174 => x"20",
   175 => x"73",
   176 => x"61",
   177 => x"6e",
   178 => x"69",
   179 => x"74",
   180 => x"79",
   181 => x"20",
   182 => x"63",
   183 => x"68",
   184 => x"65",
   185 => x"63",
   186 => x"6b",
   187 => x"2e",
   188 => x"2e",
   189 => x"2e",
   190 => x"0d",
   191 => x"0a",
   192 => x"00",
   193 => x"53",
   194 => x"61",
   195 => x"6e",
   196 => x"69",
   197 => x"74",
   198 => x"79",
   199 => x"20",
   200 => x"63",
   201 => x"68",
   202 => x"65",
   203 => x"63",
   204 => x"6b",
   205 => x"20",
   206 => x"70",
   207 => x"61",
   208 => x"73",
   209 => x"73",
   210 => x"65",
   211 => x"64",
   212 => x"2e",
   213 => x"0d",
   214 => x"0a",
   215 => x"00",
   216 => x"53",
   217 => x"61",
   218 => x"6e",
   219 => x"69",
   220 => x"74",
   221 => x"79",
   222 => x"20",
   223 => x"63",
   224 => x"68",
   225 => x"65",
   226 => x"63",
   227 => x"6b",
   228 => x"20",
   229 => x"66",
   230 => x"61",
   231 => x"69",
   232 => x"6c",
   233 => x"65",
   234 => x"64",
   235 => x"2e",
   236 => x"0d",
   237 => x"0a",
   238 => x"00",
   239 => x"00",
   240 => x"c0",
   241 => x"bc",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"df",
   246 => x"90",
   247 => x"3c",
   248 => x"00",
   249 => x"37",
   250 => x"6a",
   251 => x"04",
   252 => x"d0",
   253 => x"3c",
   254 => x"00",
   255 => x"27",
   256 => x"e9",
   257 => x"8e",
   258 => x"8c",
   259 => x"00",
   260 => x"20",
   261 => x"86",
   262 => x"4e",
   263 => x"75",
   264 => x"c0",
   265 => x"bc",
   266 => x"00",
   267 => x"00",
   268 => x"00",
   269 => x"df",
   270 => x"90",
   271 => x"3c",
   272 => x"00",
   273 => x"37",
   274 => x"6a",
   275 => x"04",
   276 => x"d0",
   277 => x"3c",
   278 => x"00",
   279 => x"27",
   280 => x"e9",
   281 => x"0f",
   282 => x"8e",
   283 => x"00",
   284 => x"10",
   285 => x"87",
   286 => x"4e",
   287 => x"75",
   288 => x"52",
   289 => x"79",
   290 => x"00",
   291 => x"7f",
   292 => x"00",
   293 => x"0c",
   294 => x"b0",
   295 => x"3c",
   296 => x"00",
   297 => x"53",
   298 => x"66",
   299 => x"2a",
   300 => x"33",
   301 => x"fc",
   302 => x"ff",
   303 => x"ff",
   304 => x"81",
   305 => x"00",
   306 => x"00",
   307 => x"06",
   308 => x"72",
   309 => x"00",
   310 => x"2e",
   311 => x"01",
   312 => x"2c",
   313 => x"01",
   314 => x"33",
   315 => x"c1",
   316 => x"00",
   317 => x"7f",
   318 => x"00",
   319 => x"0c",
   320 => x"23",
   321 => x"c1",
   322 => x"00",
   323 => x"7f",
   324 => x"00",
   325 => x"08",
   326 => x"23",
   327 => x"c1",
   328 => x"00",
   329 => x"7f",
   330 => x"00",
   331 => x"04",
   332 => x"23",
   333 => x"c1",
   334 => x"00",
   335 => x"7f",
   336 => x"00",
   337 => x"10",
   338 => x"60",
   339 => x"00",
   340 => x"01",
   341 => x"72",
   342 => x"2c",
   343 => x"39",
   344 => x"00",
   345 => x"7f",
   346 => x"00",
   347 => x"20",
   348 => x"2e",
   349 => x"39",
   350 => x"00",
   351 => x"7f",
   352 => x"00",
   353 => x"1c",
   354 => x"0c",
   355 => x"79",
   356 => x"00",
   357 => x"01",
   358 => x"00",
   359 => x"7f",
   360 => x"00",
   361 => x"0c",
   362 => x"66",
   363 => x"34",
   364 => x"33",
   365 => x"fc",
   366 => x"f0",
   367 => x"00",
   368 => x"81",
   369 => x"00",
   370 => x"00",
   371 => x"06",
   372 => x"41",
   373 => x"f9",
   374 => x"00",
   375 => x"7f",
   376 => x"00",
   377 => x"13",
   378 => x"61",
   379 => x"8c",
   380 => x"22",
   381 => x"39",
   382 => x"00",
   383 => x"7f",
   384 => x"00",
   385 => x"10",
   386 => x"b2",
   387 => x"bc",
   388 => x"00",
   389 => x"00",
   390 => x"00",
   391 => x"03",
   392 => x"6f",
   393 => x"08",
   394 => x"72",
   395 => x"0a",
   396 => x"92",
   397 => x"b9",
   398 => x"00",
   399 => x"7f",
   400 => x"00",
   401 => x"10",
   402 => x"52",
   403 => x"81",
   404 => x"e3",
   405 => x"89",
   406 => x"23",
   407 => x"c1",
   408 => x"00",
   409 => x"7f",
   410 => x"00",
   411 => x"14",
   412 => x"60",
   413 => x"00",
   414 => x"01",
   415 => x"28",
   416 => x"33",
   417 => x"f9",
   418 => x"00",
   419 => x"7f",
   420 => x"00",
   421 => x"12",
   422 => x"81",
   423 => x"00",
   424 => x"00",
   425 => x"06",
   426 => x"4a",
   427 => x"b9",
   428 => x"00",
   429 => x"7f",
   430 => x"00",
   431 => x"10",
   432 => x"67",
   433 => x"00",
   434 => x"01",
   435 => x"14",
   436 => x"0c",
   437 => x"b9",
   438 => x"00",
   439 => x"00",
   440 => x"00",
   441 => x"09",
   442 => x"00",
   443 => x"7f",
   444 => x"00",
   445 => x"10",
   446 => x"6e",
   447 => x"00",
   448 => x"00",
   449 => x"c0",
   450 => x"0c",
   451 => x"79",
   452 => x"00",
   453 => x"03",
   454 => x"00",
   455 => x"7f",
   456 => x"00",
   457 => x"0c",
   458 => x"6e",
   459 => x"16",
   460 => x"33",
   461 => x"fc",
   462 => x"0f",
   463 => x"00",
   464 => x"81",
   465 => x"00",
   466 => x"00",
   467 => x"06",
   468 => x"41",
   469 => x"f9",
   470 => x"00",
   471 => x"7f",
   472 => x"00",
   473 => x"07",
   474 => x"61",
   475 => x"00",
   476 => x"ff",
   477 => x"2c",
   478 => x"60",
   479 => x"00",
   480 => x"00",
   481 => x"e6",
   482 => x"22",
   483 => x"39",
   484 => x"00",
   485 => x"7f",
   486 => x"00",
   487 => x"14",
   488 => x"56",
   489 => x"41",
   490 => x"34",
   491 => x"39",
   492 => x"00",
   493 => x"7f",
   494 => x"00",
   495 => x"0c",
   496 => x"b4",
   497 => x"41",
   498 => x"6e",
   499 => x"20",
   500 => x"41",
   501 => x"f9",
   502 => x"00",
   503 => x"7f",
   504 => x"00",
   505 => x"08",
   506 => x"61",
   507 => x"00",
   508 => x"fe",
   509 => x"f4",
   510 => x"33",
   511 => x"f9",
   512 => x"00",
   513 => x"7f",
   514 => x"00",
   515 => x"0a",
   516 => x"81",
   517 => x"00",
   518 => x"00",
   519 => x"06",
   520 => x"33",
   521 => x"fc",
   522 => x"00",
   523 => x"01",
   524 => x"00",
   525 => x"7f",
   526 => x"00",
   527 => x"18",
   528 => x"60",
   529 => x"00",
   530 => x"00",
   531 => x"b4",
   532 => x"0c",
   533 => x"b9",
   534 => x"00",
   535 => x"00",
   536 => x"00",
   537 => x"03",
   538 => x"00",
   539 => x"7f",
   540 => x"00",
   541 => x"10",
   542 => x"6e",
   543 => x"60",
   544 => x"33",
   545 => x"fc",
   546 => x"00",
   547 => x"0f",
   548 => x"81",
   549 => x"00",
   550 => x"00",
   551 => x"06",
   552 => x"22",
   553 => x"39",
   554 => x"00",
   555 => x"7f",
   556 => x"00",
   557 => x"04",
   558 => x"e3",
   559 => x"89",
   560 => x"52",
   561 => x"81",
   562 => x"34",
   563 => x"39",
   564 => x"00",
   565 => x"7f",
   566 => x"00",
   567 => x"0c",
   568 => x"b4",
   569 => x"41",
   570 => x"6e",
   571 => x"2a",
   572 => x"20",
   573 => x"79",
   574 => x"00",
   575 => x"7f",
   576 => x"00",
   577 => x"08",
   578 => x"61",
   579 => x"00",
   580 => x"fe",
   581 => x"c4",
   582 => x"32",
   583 => x"39",
   584 => x"00",
   585 => x"7f",
   586 => x"00",
   587 => x"18",
   588 => x"53",
   589 => x"79",
   590 => x"00",
   591 => x"7f",
   592 => x"00",
   593 => x"18",
   594 => x"53",
   595 => x"41",
   596 => x"6a",
   597 => x"70",
   598 => x"52",
   599 => x"b9",
   600 => x"00",
   601 => x"7f",
   602 => x"00",
   603 => x"08",
   604 => x"33",
   605 => x"fc",
   606 => x"00",
   607 => x"01",
   608 => x"00",
   609 => x"7f",
   610 => x"00",
   611 => x"18",
   612 => x"60",
   613 => x"60",
   614 => x"30",
   615 => x"39",
   616 => x"00",
   617 => x"7f",
   618 => x"00",
   619 => x"18",
   620 => x"52",
   621 => x"40",
   622 => x"c0",
   623 => x"7c",
   624 => x"00",
   625 => x"01",
   626 => x"67",
   627 => x"52",
   628 => x"20",
   629 => x"79",
   630 => x"00",
   631 => x"7f",
   632 => x"00",
   633 => x"08",
   634 => x"e5",
   635 => x"88",
   636 => x"e1",
   637 => x"2f",
   638 => x"10",
   639 => x"87",
   640 => x"33",
   641 => x"fc",
   642 => x"f0",
   643 => x"f0",
   644 => x"81",
   645 => x"00",
   646 => x"00",
   647 => x"06",
   648 => x"0c",
   649 => x"b9",
   650 => x"00",
   651 => x"00",
   652 => x"00",
   653 => x"07",
   654 => x"00",
   655 => x"7f",
   656 => x"00",
   657 => x"10",
   658 => x"6d",
   659 => x"32",
   660 => x"33",
   661 => x"fc",
   662 => x"f0",
   663 => x"0f",
   664 => x"81",
   665 => x"00",
   666 => x"00",
   667 => x"06",
   668 => x"0c",
   669 => x"b9",
   670 => x"00",
   671 => x"00",
   672 => x"00",
   673 => x"09",
   674 => x"00",
   675 => x"7f",
   676 => x"00",
   677 => x"10",
   678 => x"6e",
   679 => x"1e",
   680 => x"33",
   681 => x"fc",
   682 => x"ff",
   683 => x"f0",
   684 => x"81",
   685 => x"00",
   686 => x"00",
   687 => x"06",
   688 => x"41",
   689 => x"fa",
   690 => x"00",
   691 => x"22",
   692 => x"61",
   693 => x"56",
   694 => x"2e",
   695 => x"b9",
   696 => x"00",
   697 => x"7f",
   698 => x"00",
   699 => x"08",
   700 => x"08",
   701 => x"b9",
   702 => x"00",
   703 => x"00",
   704 => x"81",
   705 => x"00",
   706 => x"00",
   707 => x"04",
   708 => x"4e",
   709 => x"75",
   710 => x"23",
   711 => x"c6",
   712 => x"00",
   713 => x"7f",
   714 => x"00",
   715 => x"20",
   716 => x"23",
   717 => x"c7",
   718 => x"00",
   719 => x"7f",
   720 => x"00",
   721 => x"1c",
   722 => x"4e",
   723 => x"75",
   724 => x"46",
   725 => x"69",
   726 => x"72",
   727 => x"6d",
   728 => x"77",
   729 => x"61",
   730 => x"72",
   731 => x"65",
   732 => x"20",
   733 => x"72",
   734 => x"65",
   735 => x"63",
   736 => x"65",
   737 => x"69",
   738 => x"76",
   739 => x"65",
   740 => x"64",
   741 => x"20",
   742 => x"2d",
   743 => x"20",
   744 => x"6c",
   745 => x"61",
   746 => x"75",
   747 => x"6e",
   748 => x"63",
   749 => x"68",
   750 => x"69",
   751 => x"6e",
   752 => x"67",
   753 => x"0d",
   754 => x"0a",
   755 => x"00",
   756 => x"48",
   757 => x"40",
   758 => x"30",
   759 => x"39",
   760 => x"81",
   761 => x"00",
   762 => x"00",
   763 => x"00",
   764 => x"08",
   765 => x"00",
   766 => x"00",
   767 => x"08",
   768 => x"67",
   769 => x"f4",
   770 => x"48",
   771 => x"40",
   772 => x"33",
   773 => x"c0",
   774 => x"81",
   775 => x"00",
   776 => x"00",
   777 => x"00",
   778 => x"4e",
   779 => x"75",
   780 => x"2f",
   781 => x"00",
   782 => x"70",
   783 => x"00",
   784 => x"30",
   785 => x"39",
   786 => x"81",
   787 => x"00",
   788 => x"00",
   789 => x"00",
   790 => x"08",
   791 => x"00",
   792 => x"00",
   793 => x"08",
   794 => x"67",
   795 => x"f4",
   796 => x"10",
   797 => x"18",
   798 => x"67",
   799 => x"08",
   800 => x"33",
   801 => x"c0",
   802 => x"81",
   803 => x"00",
   804 => x"00",
   805 => x"00",
   806 => x"60",
   807 => x"e8",
   808 => x"20",
   809 => x"1f",
   810 => x"4e",
   811 => x"75",
   812 => x"33",
   813 => x"fc",
   814 => x"00",
   815 => x"01",
   816 => x"81",
   817 => x"00",
   818 => x"00",
   819 => x"06",
   820 => x"41",
   821 => x"fa",
   822 => x"01",
   823 => x"fa",
   824 => x"61",
   825 => x"00",
   826 => x"03",
   827 => x"e2",
   828 => x"61",
   829 => x"00",
   830 => x"02",
   831 => x"60",
   832 => x"66",
   833 => x"5c",
   834 => x"33",
   835 => x"fc",
   836 => x"00",
   837 => x"02",
   838 => x"81",
   839 => x"00",
   840 => x"00",
   841 => x"06",
   842 => x"33",
   843 => x"fc",
   844 => x"00",
   845 => x"40",
   846 => x"00",
   847 => x"7f",
   848 => x"00",
   849 => x"26",
   850 => x"61",
   851 => x"00",
   852 => x"04",
   853 => x"8a",
   854 => x"67",
   855 => x"0c",
   856 => x"42",
   857 => x"79",
   858 => x"00",
   859 => x"7f",
   860 => x"00",
   861 => x"26",
   862 => x"61",
   863 => x"00",
   864 => x"04",
   865 => x"7e",
   866 => x"66",
   867 => x"28",
   868 => x"33",
   869 => x"fc",
   870 => x"00",
   871 => x"03",
   872 => x"81",
   873 => x"00",
   874 => x"00",
   875 => x"06",
   876 => x"61",
   877 => x"00",
   878 => x"05",
   879 => x"f8",
   880 => x"43",
   881 => x"fa",
   882 => x"00",
   883 => x"57",
   884 => x"61",
   885 => x"00",
   886 => x"06",
   887 => x"48",
   888 => x"67",
   889 => x"12",
   890 => x"41",
   891 => x"fa",
   892 => x"00",
   893 => x"47",
   894 => x"61",
   895 => x"00",
   896 => x"03",
   897 => x"9c",
   898 => x"30",
   899 => x"7c",
   900 => x"20",
   901 => x"00",
   902 => x"61",
   903 => x"00",
   904 => x"04",
   905 => x"02",
   906 => x"4e",
   907 => x"75",
   908 => x"33",
   909 => x"fc",
   910 => x"f0",
   911 => x"03",
   912 => x"81",
   913 => x"00",
   914 => x"00",
   915 => x"06",
   916 => x"41",
   917 => x"fa",
   918 => x"00",
   919 => x"29",
   920 => x"61",
   921 => x"00",
   922 => x"03",
   923 => x"82",
   924 => x"4e",
   925 => x"75",
   926 => x"33",
   927 => x"fc",
   928 => x"f0",
   929 => x"02",
   930 => x"81",
   931 => x"00",
   932 => x"00",
   933 => x"06",
   934 => x"41",
   935 => x"fa",
   936 => x"00",
   937 => x"08",
   938 => x"61",
   939 => x"00",
   940 => x"03",
   941 => x"70",
   942 => x"4e",
   943 => x"75",
   944 => x"53",
   945 => x"44",
   946 => x"20",
   947 => x"69",
   948 => x"6e",
   949 => x"69",
   950 => x"74",
   951 => x"20",
   952 => x"66",
   953 => x"61",
   954 => x"69",
   955 => x"6c",
   956 => x"65",
   957 => x"64",
   958 => x"00",
   959 => x"6e",
   960 => x"6f",
   961 => x"74",
   962 => x"20",
   963 => x"66",
   964 => x"6f",
   965 => x"75",
   966 => x"6e",
   967 => x"64",
   968 => x"20",
   969 => x"42",
   970 => x"4f",
   971 => x"4f",
   972 => x"54",
   973 => x"20",
   974 => x"20",
   975 => x"20",
   976 => x"20",
   977 => x"53",
   978 => x"52",
   979 => x"45",
   980 => x"00",
   981 => x"00",
   982 => x"33",
   983 => x"fc",
   984 => x"01",
   985 => x"00",
   986 => x"81",
   987 => x"00",
   988 => x"00",
   989 => x"06",
   990 => x"41",
   991 => x"f9",
   992 => x"00",
   993 => x"7f",
   994 => x"00",
   995 => x"56",
   996 => x"61",
   997 => x"00",
   998 => x"00",
   999 => x"c4",
  1000 => x"66",
  1001 => x"68",
  1002 => x"33",
  1003 => x"fc",
  1004 => x"01",
  1005 => x"01",
  1006 => x"81",
  1007 => x"00",
  1008 => x"00",
  1009 => x"06",
  1010 => x"32",
  1011 => x"3c",
  1012 => x"4e",
  1013 => x"20",
  1014 => x"53",
  1015 => x"41",
  1016 => x"67",
  1017 => x"44",
  1018 => x"33",
  1019 => x"fc",
  1020 => x"01",
  1021 => x"02",
  1022 => x"81",
  1023 => x"00",
  1024 => x"00",
  1025 => x"06",
  1026 => x"33",
  1027 => x"7c",
  1028 => x"00",
  1029 => x"ff",
  1030 => x"00",
  1031 => x"24",
  1032 => x"30",
  1033 => x"29",
  1034 => x"00",
  1035 => x"24",
  1036 => x"b0",
  1037 => x"3c",
  1038 => x"00",
  1039 => x"fe",
  1040 => x"66",
  1041 => x"e4",
  1042 => x"30",
  1043 => x"29",
  1044 => x"01",
  1045 => x"00",
  1046 => x"32",
  1047 => x"3c",
  1048 => x"00",
  1049 => x"7f",
  1050 => x"20",
  1051 => x"29",
  1052 => x"01",
  1053 => x"00",
  1054 => x"20",
  1055 => x"c0",
  1056 => x"51",
  1057 => x"c9",
  1058 => x"ff",
  1059 => x"f8",
  1060 => x"30",
  1061 => x"29",
  1062 => x"00",
  1063 => x"24",
  1064 => x"33",
  1065 => x"7c",
  1066 => x"00",
  1067 => x"00",
  1068 => x"00",
  1069 => x"22",
  1070 => x"33",
  1071 => x"fc",
  1072 => x"01",
  1073 => x"03",
  1074 => x"81",
  1075 => x"00",
  1076 => x"00",
  1077 => x"06",
  1078 => x"41",
  1079 => x"e8",
  1080 => x"fe",
  1081 => x"00",
  1082 => x"70",
  1083 => x"00",
  1084 => x"4e",
  1085 => x"75",
  1086 => x"33",
  1087 => x"fc",
  1088 => x"f1",
  1089 => x"02",
  1090 => x"81",
  1091 => x"00",
  1092 => x"00",
  1093 => x"06",
  1094 => x"41",
  1095 => x"fa",
  1096 => x"01",
  1097 => x"38",
  1098 => x"61",
  1099 => x"00",
  1100 => x"02",
  1101 => x"d0",
  1102 => x"70",
  1103 => x"fe",
  1104 => x"4e",
  1105 => x"75",
  1106 => x"33",
  1107 => x"fc",
  1108 => x"f1",
  1109 => x"03",
  1110 => x"81",
  1111 => x"00",
  1112 => x"00",
  1113 => x"06",
  1114 => x"41",
  1115 => x"fa",
  1116 => x"01",
  1117 => x"0c",
  1118 => x"61",
  1119 => x"00",
  1120 => x"02",
  1121 => x"bc",
  1122 => x"70",
  1123 => x"ff",
  1124 => x"4e",
  1125 => x"75",
  1126 => x"22",
  1127 => x"3c",
  1128 => x"00",
  1129 => x"95",
  1130 => x"00",
  1131 => x"40",
  1132 => x"70",
  1133 => x"00",
  1134 => x"60",
  1135 => x"40",
  1136 => x"22",
  1137 => x"3c",
  1138 => x"00",
  1139 => x"ff",
  1140 => x"00",
  1141 => x"41",
  1142 => x"70",
  1143 => x"00",
  1144 => x"60",
  1145 => x"36",
  1146 => x"22",
  1147 => x"3c",
  1148 => x"00",
  1149 => x"87",
  1150 => x"00",
  1151 => x"48",
  1152 => x"20",
  1153 => x"3c",
  1154 => x"00",
  1155 => x"00",
  1156 => x"01",
  1157 => x"aa",
  1158 => x"60",
  1159 => x"28",
  1160 => x"22",
  1161 => x"3c",
  1162 => x"00",
  1163 => x"87",
  1164 => x"00",
  1165 => x"69",
  1166 => x"20",
  1167 => x"3c",
  1168 => x"40",
  1169 => x"00",
  1170 => x"00",
  1171 => x"00",
  1172 => x"60",
  1173 => x"1a",
  1174 => x"22",
  1175 => x"3c",
  1176 => x"00",
  1177 => x"ff",
  1178 => x"00",
  1179 => x"77",
  1180 => x"70",
  1181 => x"00",
  1182 => x"60",
  1183 => x"10",
  1184 => x"22",
  1185 => x"3c",
  1186 => x"00",
  1187 => x"ff",
  1188 => x"00",
  1189 => x"7a",
  1190 => x"70",
  1191 => x"00",
  1192 => x"60",
  1193 => x"06",
  1194 => x"22",
  1195 => x"3c",
  1196 => x"00",
  1197 => x"ff",
  1198 => x"00",
  1199 => x"51",
  1200 => x"43",
  1201 => x"f9",
  1202 => x"81",
  1203 => x"00",
  1204 => x"00",
  1205 => x"00",
  1206 => x"33",
  1207 => x"7c",
  1208 => x"00",
  1209 => x"ff",
  1210 => x"00",
  1211 => x"24",
  1212 => x"3f",
  1213 => x"69",
  1214 => x"00",
  1215 => x"24",
  1216 => x"ff",
  1217 => x"fe",
  1218 => x"33",
  1219 => x"7c",
  1220 => x"00",
  1221 => x"01",
  1222 => x"00",
  1223 => x"22",
  1224 => x"33",
  1225 => x"7c",
  1226 => x"00",
  1227 => x"ff",
  1228 => x"00",
  1229 => x"24",
  1230 => x"33",
  1231 => x"41",
  1232 => x"00",
  1233 => x"24",
  1234 => x"48",
  1235 => x"41",
  1236 => x"4a",
  1237 => x"79",
  1238 => x"00",
  1239 => x"7f",
  1240 => x"00",
  1241 => x"24",
  1242 => x"67",
  1243 => x"16",
  1244 => x"e1",
  1245 => x"98",
  1246 => x"33",
  1247 => x"40",
  1248 => x"00",
  1249 => x"24",
  1250 => x"e1",
  1251 => x"98",
  1252 => x"33",
  1253 => x"40",
  1254 => x"00",
  1255 => x"24",
  1256 => x"e1",
  1257 => x"98",
  1258 => x"33",
  1259 => x"40",
  1260 => x"00",
  1261 => x"24",
  1262 => x"e1",
  1263 => x"98",
  1264 => x"60",
  1265 => x"18",
  1266 => x"d0",
  1267 => x"80",
  1268 => x"48",
  1269 => x"40",
  1270 => x"33",
  1271 => x"40",
  1272 => x"00",
  1273 => x"24",
  1274 => x"48",
  1275 => x"40",
  1276 => x"e1",
  1277 => x"58",
  1278 => x"33",
  1279 => x"40",
  1280 => x"00",
  1281 => x"24",
  1282 => x"e1",
  1283 => x"58",
  1284 => x"33",
  1285 => x"40",
  1286 => x"00",
  1287 => x"24",
  1288 => x"70",
  1289 => x"00",
  1290 => x"33",
  1291 => x"40",
  1292 => x"00",
  1293 => x"24",
  1294 => x"33",
  1295 => x"41",
  1296 => x"00",
  1297 => x"24",
  1298 => x"22",
  1299 => x"3c",
  1300 => x"00",
  1301 => x"00",
  1302 => x"01",
  1303 => x"90",
  1304 => x"53",
  1305 => x"81",
  1306 => x"67",
  1307 => x"10",
  1308 => x"33",
  1309 => x"7c",
  1310 => x"00",
  1311 => x"ff",
  1312 => x"00",
  1313 => x"24",
  1314 => x"30",
  1315 => x"29",
  1316 => x"00",
  1317 => x"24",
  1318 => x"b0",
  1319 => x"3c",
  1320 => x"00",
  1321 => x"ff",
  1322 => x"67",
  1323 => x"ec",
  1324 => x"80",
  1325 => x"00",
  1326 => x"4e",
  1327 => x"75",
  1328 => x"53",
  1329 => x"74",
  1330 => x"61",
  1331 => x"72",
  1332 => x"74",
  1333 => x"20",
  1334 => x"49",
  1335 => x"6e",
  1336 => x"69",
  1337 => x"74",
  1338 => x"0d",
  1339 => x"0a",
  1340 => x"00",
  1341 => x"49",
  1342 => x"6e",
  1343 => x"69",
  1344 => x"74",
  1345 => x"20",
  1346 => x"64",
  1347 => x"6f",
  1348 => x"6e",
  1349 => x"65",
  1350 => x"0d",
  1351 => x"0a",
  1352 => x"00",
  1353 => x"49",
  1354 => x"6e",
  1355 => x"69",
  1356 => x"74",
  1357 => x"20",
  1358 => x"66",
  1359 => x"61",
  1360 => x"69",
  1361 => x"6c",
  1362 => x"75",
  1363 => x"72",
  1364 => x"65",
  1365 => x"0d",
  1366 => x"0a",
  1367 => x"00",
  1368 => x"52",
  1369 => x"65",
  1370 => x"73",
  1371 => x"65",
  1372 => x"74",
  1373 => x"20",
  1374 => x"66",
  1375 => x"61",
  1376 => x"69",
  1377 => x"6c",
  1378 => x"75",
  1379 => x"72",
  1380 => x"65",
  1381 => x"0d",
  1382 => x"0a",
  1383 => x"00",
  1384 => x"43",
  1385 => x"6f",
  1386 => x"6d",
  1387 => x"6d",
  1388 => x"61",
  1389 => x"6e",
  1390 => x"64",
  1391 => x"20",
  1392 => x"54",
  1393 => x"69",
  1394 => x"6d",
  1395 => x"65",
  1396 => x"6f",
  1397 => x"75",
  1398 => x"74",
  1399 => x"5f",
  1400 => x"45",
  1401 => x"72",
  1402 => x"72",
  1403 => x"6f",
  1404 => x"72",
  1405 => x"0d",
  1406 => x"0a",
  1407 => x"00",
  1408 => x"54",
  1409 => x"69",
  1410 => x"6d",
  1411 => x"65",
  1412 => x"6f",
  1413 => x"75",
  1414 => x"74",
  1415 => x"5f",
  1416 => x"45",
  1417 => x"72",
  1418 => x"72",
  1419 => x"6f",
  1420 => x"72",
  1421 => x"0d",
  1422 => x"0a",
  1423 => x"00",
  1424 => x"53",
  1425 => x"44",
  1426 => x"48",
  1427 => x"43",
  1428 => x"20",
  1429 => x"66",
  1430 => x"6f",
  1431 => x"75",
  1432 => x"6e",
  1433 => x"64",
  1434 => x"20",
  1435 => x"0d",
  1436 => x"0a",
  1437 => x"00",
  1438 => x"33",
  1439 => x"fc",
  1440 => x"ff",
  1441 => x"ff",
  1442 => x"00",
  1443 => x"7f",
  1444 => x"00",
  1445 => x"24",
  1446 => x"43",
  1447 => x"f9",
  1448 => x"81",
  1449 => x"00",
  1450 => x"00",
  1451 => x"00",
  1452 => x"33",
  1453 => x"7c",
  1454 => x"00",
  1455 => x"00",
  1456 => x"00",
  1457 => x"22",
  1458 => x"33",
  1459 => x"7c",
  1460 => x"00",
  1461 => x"96",
  1462 => x"00",
  1463 => x"1e",
  1464 => x"32",
  1465 => x"3c",
  1466 => x"00",
  1467 => x"c8",
  1468 => x"43",
  1469 => x"e9",
  1470 => x"00",
  1471 => x"20",
  1472 => x"33",
  1473 => x"7c",
  1474 => x"00",
  1475 => x"ff",
  1476 => x"00",
  1477 => x"24",
  1478 => x"51",
  1479 => x"c9",
  1480 => x"ff",
  1481 => x"f8",
  1482 => x"34",
  1483 => x"3c",
  1484 => x"00",
  1485 => x"32",
  1486 => x"61",
  1487 => x"00",
  1488 => x"fe",
  1489 => x"96",
  1490 => x"3f",
  1491 => x"69",
  1492 => x"00",
  1493 => x"24",
  1494 => x"ff",
  1495 => x"fe",
  1496 => x"33",
  1497 => x"7c",
  1498 => x"00",
  1499 => x"00",
  1500 => x"00",
  1501 => x"22",
  1502 => x"b0",
  1503 => x"3c",
  1504 => x"00",
  1505 => x"01",
  1506 => x"67",
  1507 => x"12",
  1508 => x"51",
  1509 => x"ca",
  1510 => x"ff",
  1511 => x"e8",
  1512 => x"48",
  1513 => x"7a",
  1514 => x"ff",
  1515 => x"6e",
  1516 => x"61",
  1517 => x"00",
  1518 => x"01",
  1519 => x"22",
  1520 => x"58",
  1521 => x"8f",
  1522 => x"70",
  1523 => x"ff",
  1524 => x"4e",
  1525 => x"75",
  1526 => x"22",
  1527 => x"3c",
  1528 => x"00",
  1529 => x"00",
  1530 => x"20",
  1531 => x"00",
  1532 => x"33",
  1533 => x"7c",
  1534 => x"00",
  1535 => x"ff",
  1536 => x"00",
  1537 => x"24",
  1538 => x"53",
  1539 => x"81",
  1540 => x"66",
  1541 => x"f6",
  1542 => x"61",
  1543 => x"00",
  1544 => x"fe",
  1545 => x"72",
  1546 => x"b0",
  1547 => x"3c",
  1548 => x"00",
  1549 => x"01",
  1550 => x"66",
  1551 => x"00",
  1552 => x"00",
  1553 => x"9e",
  1554 => x"33",
  1555 => x"7c",
  1556 => x"00",
  1557 => x"ff",
  1558 => x"00",
  1559 => x"24",
  1560 => x"33",
  1561 => x"7c",
  1562 => x"00",
  1563 => x"ff",
  1564 => x"00",
  1565 => x"24",
  1566 => x"33",
  1567 => x"7c",
  1568 => x"00",
  1569 => x"ff",
  1570 => x"00",
  1571 => x"24",
  1572 => x"30",
  1573 => x"29",
  1574 => x"00",
  1575 => x"24",
  1576 => x"0c",
  1577 => x"00",
  1578 => x"00",
  1579 => x"01",
  1580 => x"66",
  1581 => x"00",
  1582 => x"00",
  1583 => x"80",
  1584 => x"33",
  1585 => x"7c",
  1586 => x"00",
  1587 => x"ff",
  1588 => x"00",
  1589 => x"24",
  1590 => x"30",
  1591 => x"29",
  1592 => x"00",
  1593 => x"24",
  1594 => x"0c",
  1595 => x"00",
  1596 => x"00",
  1597 => x"aa",
  1598 => x"66",
  1599 => x"6e",
  1600 => x"3f",
  1601 => x"69",
  1602 => x"00",
  1603 => x"24",
  1604 => x"ff",
  1605 => x"fe",
  1606 => x"33",
  1607 => x"7c",
  1608 => x"00",
  1609 => x"00",
  1610 => x"00",
  1611 => x"22",
  1612 => x"48",
  1613 => x"7a",
  1614 => x"ff",
  1615 => x"42",
  1616 => x"61",
  1617 => x"00",
  1618 => x"00",
  1619 => x"be",
  1620 => x"58",
  1621 => x"8f",
  1622 => x"34",
  1623 => x"3c",
  1624 => x"00",
  1625 => x"32",
  1626 => x"53",
  1627 => x"42",
  1628 => x"67",
  1629 => x"50",
  1630 => x"32",
  1631 => x"3c",
  1632 => x"07",
  1633 => x"d0",
  1634 => x"33",
  1635 => x"7c",
  1636 => x"00",
  1637 => x"ff",
  1638 => x"00",
  1639 => x"24",
  1640 => x"51",
  1641 => x"c9",
  1642 => x"ff",
  1643 => x"f8",
  1644 => x"61",
  1645 => x"00",
  1646 => x"fe",
  1647 => x"28",
  1648 => x"b0",
  1649 => x"3c",
  1650 => x"00",
  1651 => x"01",
  1652 => x"66",
  1653 => x"e4",
  1654 => x"61",
  1655 => x"00",
  1656 => x"fe",
  1657 => x"10",
  1658 => x"66",
  1659 => x"de",
  1660 => x"61",
  1661 => x"00",
  1662 => x"fe",
  1663 => x"22",
  1664 => x"66",
  1665 => x"d8",
  1666 => x"33",
  1667 => x"7c",
  1668 => x"00",
  1669 => x"ff",
  1670 => x"00",
  1671 => x"24",
  1672 => x"30",
  1673 => x"29",
  1674 => x"00",
  1675 => x"24",
  1676 => x"c0",
  1677 => x"3c",
  1678 => x"00",
  1679 => x"40",
  1680 => x"66",
  1681 => x"08",
  1682 => x"33",
  1683 => x"fc",
  1684 => x"00",
  1685 => x"00",
  1686 => x"00",
  1687 => x"7f",
  1688 => x"00",
  1689 => x"24",
  1690 => x"33",
  1691 => x"7c",
  1692 => x"00",
  1693 => x"ff",
  1694 => x"00",
  1695 => x"24",
  1696 => x"33",
  1697 => x"7c",
  1698 => x"00",
  1699 => x"ff",
  1700 => x"00",
  1701 => x"24",
  1702 => x"33",
  1703 => x"7c",
  1704 => x"00",
  1705 => x"ff",
  1706 => x"00",
  1707 => x"24",
  1708 => x"60",
  1709 => x"3c",
  1710 => x"33",
  1711 => x"fc",
  1712 => x"00",
  1713 => x"00",
  1714 => x"00",
  1715 => x"7f",
  1716 => x"00",
  1717 => x"24",
  1718 => x"34",
  1719 => x"3c",
  1720 => x"00",
  1721 => x"0a",
  1722 => x"32",
  1723 => x"3c",
  1724 => x"07",
  1725 => x"d0",
  1726 => x"33",
  1727 => x"7c",
  1728 => x"00",
  1729 => x"ff",
  1730 => x"00",
  1731 => x"24",
  1732 => x"51",
  1733 => x"c9",
  1734 => x"ff",
  1735 => x"f8",
  1736 => x"61",
  1737 => x"00",
  1738 => x"fd",
  1739 => x"a6",
  1740 => x"67",
  1741 => x"1c",
  1742 => x"3f",
  1743 => x"69",
  1744 => x"00",
  1745 => x"24",
  1746 => x"ff",
  1747 => x"fe",
  1748 => x"33",
  1749 => x"7c",
  1750 => x"00",
  1751 => x"00",
  1752 => x"00",
  1753 => x"22",
  1754 => x"51",
  1755 => x"ca",
  1756 => x"ff",
  1757 => x"de",
  1758 => x"48",
  1759 => x"7a",
  1760 => x"fe",
  1761 => x"69",
  1762 => x"61",
  1763 => x"2c",
  1764 => x"58",
  1765 => x"8f",
  1766 => x"70",
  1767 => x"ff",
  1768 => x"4e",
  1769 => x"75",
  1770 => x"3f",
  1771 => x"69",
  1772 => x"00",
  1773 => x"24",
  1774 => x"ff",
  1775 => x"fe",
  1776 => x"33",
  1777 => x"7c",
  1778 => x"00",
  1779 => x"00",
  1780 => x"00",
  1781 => x"22",
  1782 => x"33",
  1783 => x"69",
  1784 => x"00",
  1785 => x"2c",
  1786 => x"00",
  1787 => x"1e",
  1788 => x"48",
  1789 => x"7a",
  1790 => x"fe",
  1791 => x"3f",
  1792 => x"61",
  1793 => x"0e",
  1794 => x"58",
  1795 => x"8f",
  1796 => x"33",
  1797 => x"fc",
  1798 => x"ff",
  1799 => x"ff",
  1800 => x"81",
  1801 => x"00",
  1802 => x"00",
  1803 => x"06",
  1804 => x"70",
  1805 => x"00",
  1806 => x"4e",
  1807 => x"75",
  1808 => x"2f",
  1809 => x"08",
  1810 => x"20",
  1811 => x"6f",
  1812 => x"00",
  1813 => x"08",
  1814 => x"61",
  1815 => x"04",
  1816 => x"20",
  1817 => x"5f",
  1818 => x"4e",
  1819 => x"75",
  1820 => x"48",
  1821 => x"e7",
  1822 => x"00",
  1823 => x"c0",
  1824 => x"22",
  1825 => x"39",
  1826 => x"00",
  1827 => x"7f",
  1828 => x"00",
  1829 => x"52",
  1830 => x"43",
  1831 => x"f9",
  1832 => x"80",
  1833 => x"00",
  1834 => x"08",
  1835 => x"00",
  1836 => x"10",
  1837 => x"18",
  1838 => x"67",
  1839 => x"08",
  1840 => x"13",
  1841 => x"80",
  1842 => x"10",
  1843 => x"00",
  1844 => x"52",
  1845 => x"41",
  1846 => x"60",
  1847 => x"f4",
  1848 => x"06",
  1849 => x"b9",
  1850 => x"00",
  1851 => x"00",
  1852 => x"00",
  1853 => x"4c",
  1854 => x"00",
  1855 => x"7f",
  1856 => x"00",
  1857 => x"52",
  1858 => x"4c",
  1859 => x"df",
  1860 => x"03",
  1861 => x"00",
  1862 => x"4e",
  1863 => x"75",
  1864 => x"4a",
  1865 => x"79",
  1866 => x"00",
  1867 => x"7f",
  1868 => x"00",
  1869 => x"24",
  1870 => x"67",
  1871 => x"1e",
  1872 => x"41",
  1873 => x"fa",
  1874 => x"00",
  1875 => x"08",
  1876 => x"48",
  1877 => x"7a",
  1878 => x"00",
  1879 => x"34",
  1880 => x"60",
  1881 => x"c2",
  1882 => x"53",
  1883 => x"44",
  1884 => x"48",
  1885 => x"43",
  1886 => x"20",
  1887 => x"66",
  1888 => x"6c",
  1889 => x"61",
  1890 => x"67",
  1891 => x"20",
  1892 => x"73",
  1893 => x"74",
  1894 => x"69",
  1895 => x"6c",
  1896 => x"6c",
  1897 => x"20",
  1898 => x"73",
  1899 => x"65",
  1900 => x"74",
  1901 => x"00",
  1902 => x"41",
  1903 => x"fa",
  1904 => x"00",
  1905 => x"08",
  1906 => x"48",
  1907 => x"7a",
  1908 => x"00",
  1909 => x"16",
  1910 => x"60",
  1911 => x"a4",
  1912 => x"53",
  1913 => x"44",
  1914 => x"48",
  1915 => x"43",
  1916 => x"20",
  1917 => x"66",
  1918 => x"6c",
  1919 => x"61",
  1920 => x"67",
  1921 => x"20",
  1922 => x"63",
  1923 => x"6c",
  1924 => x"65",
  1925 => x"61",
  1926 => x"72",
  1927 => x"65",
  1928 => x"64",
  1929 => x"00",
  1930 => x"61",
  1931 => x"00",
  1932 => x"02",
  1933 => x"0a",
  1934 => x"61",
  1935 => x"00",
  1936 => x"fc",
  1937 => x"46",
  1938 => x"66",
  1939 => x"46",
  1940 => x"2e",
  1941 => x"3c",
  1942 => x"00",
  1943 => x"00",
  1944 => x"01",
  1945 => x"ff",
  1946 => x"41",
  1947 => x"f9",
  1948 => x"00",
  1949 => x"7f",
  1950 => x"00",
  1951 => x"56",
  1952 => x"43",
  1953 => x"f9",
  1954 => x"80",
  1955 => x"00",
  1956 => x"08",
  1957 => x"00",
  1958 => x"10",
  1959 => x"18",
  1960 => x"12",
  1961 => x"c0",
  1962 => x"48",
  1963 => x"e7",
  1964 => x"01",
  1965 => x"c0",
  1966 => x"61",
  1967 => x"00",
  1968 => x"f9",
  1969 => x"70",
  1970 => x"4c",
  1971 => x"df",
  1972 => x"03",
  1973 => x"80",
  1974 => x"51",
  1975 => x"cf",
  1976 => x"ff",
  1977 => x"ee",
  1978 => x"20",
  1979 => x"39",
  1980 => x"00",
  1981 => x"7f",
  1982 => x"00",
  1983 => x"38",
  1984 => x"52",
  1985 => x"80",
  1986 => x"23",
  1987 => x"c0",
  1988 => x"00",
  1989 => x"7f",
  1990 => x"00",
  1991 => x"38",
  1992 => x"53",
  1993 => x"79",
  1994 => x"00",
  1995 => x"7f",
  1996 => x"00",
  1997 => x"36",
  1998 => x"66",
  1999 => x"be",
  2000 => x"61",
  2001 => x"00",
  2002 => x"02",
  2003 => x"7a",
  2004 => x"66",
  2005 => x"b4",
  2006 => x"20",
  2007 => x"08",
  2008 => x"4e",
  2009 => x"75",
  2010 => x"70",
  2011 => x"00",
  2012 => x"4e",
  2013 => x"75",
  2014 => x"33",
  2015 => x"fc",
  2016 => x"02",
  2017 => x"01",
  2018 => x"81",
  2019 => x"00",
  2020 => x"00",
  2021 => x"06",
  2022 => x"70",
  2023 => x"00",
  2024 => x"23",
  2025 => x"c0",
  2026 => x"00",
  2027 => x"7f",
  2028 => x"00",
  2029 => x"3e",
  2030 => x"33",
  2031 => x"fc",
  2032 => x"02",
  2033 => x"11",
  2034 => x"81",
  2035 => x"00",
  2036 => x"00",
  2037 => x"06",
  2038 => x"61",
  2039 => x"00",
  2040 => x"fb",
  2041 => x"de",
  2042 => x"66",
  2043 => x"5c",
  2044 => x"33",
  2045 => x"fc",
  2046 => x"02",
  2047 => x"02",
  2048 => x"81",
  2049 => x"00",
  2050 => x"00",
  2051 => x"06",
  2052 => x"0c",
  2053 => x"28",
  2054 => x"00",
  2055 => x"55",
  2056 => x"01",
  2057 => x"fe",
  2058 => x"66",
  2059 => x"4c",
  2060 => x"0c",
  2061 => x"28",
  2062 => x"00",
  2063 => x"aa",
  2064 => x"01",
  2065 => x"ff",
  2066 => x"66",
  2067 => x"44",
  2068 => x"30",
  2069 => x"39",
  2070 => x"00",
  2071 => x"7f",
  2072 => x"00",
  2073 => x"26",
  2074 => x"c0",
  2075 => x"7c",
  2076 => x"00",
  2077 => x"70",
  2078 => x"b0",
  2079 => x"7c",
  2080 => x"00",
  2081 => x"40",
  2082 => x"64",
  2083 => x"40",
  2084 => x"43",
  2085 => x"e8",
  2086 => x"01",
  2087 => x"be",
  2088 => x"d2",
  2089 => x"c0",
  2090 => x"33",
  2091 => x"fc",
  2092 => x"02",
  2093 => x"03",
  2094 => x"81",
  2095 => x"00",
  2096 => x"00",
  2097 => x"06",
  2098 => x"20",
  2099 => x"29",
  2100 => x"00",
  2101 => x"08",
  2102 => x"e0",
  2103 => x"58",
  2104 => x"48",
  2105 => x"40",
  2106 => x"e0",
  2107 => x"58",
  2108 => x"23",
  2109 => x"c0",
  2110 => x"00",
  2111 => x"7f",
  2112 => x"00",
  2113 => x"3e",
  2114 => x"61",
  2115 => x"00",
  2116 => x"fb",
  2117 => x"92",
  2118 => x"66",
  2119 => x"10",
  2120 => x"0c",
  2121 => x"28",
  2122 => x"00",
  2123 => x"55",
  2124 => x"01",
  2125 => x"fe",
  2126 => x"66",
  2127 => x"08",
  2128 => x"0c",
  2129 => x"28",
  2130 => x"00",
  2131 => x"aa",
  2132 => x"01",
  2133 => x"ff",
  2134 => x"67",
  2135 => x"0c",
  2136 => x"33",
  2137 => x"fc",
  2138 => x"f2",
  2139 => x"01",
  2140 => x"81",
  2141 => x"00",
  2142 => x"00",
  2143 => x"06",
  2144 => x"70",
  2145 => x"ff",
  2146 => x"4e",
  2147 => x"75",
  2148 => x"33",
  2149 => x"fc",
  2150 => x"02",
  2151 => x"04",
  2152 => x"81",
  2153 => x"00",
  2154 => x"00",
  2155 => x"06",
  2156 => x"0c",
  2157 => x"a8",
  2158 => x"46",
  2159 => x"41",
  2160 => x"54",
  2161 => x"31",
  2162 => x"00",
  2163 => x"36",
  2164 => x"66",
  2165 => x"24",
  2166 => x"13",
  2167 => x"fc",
  2168 => x"00",
  2169 => x"0c",
  2170 => x"00",
  2171 => x"7f",
  2172 => x"00",
  2173 => x"28",
  2174 => x"0c",
  2175 => x"a8",
  2176 => x"32",
  2177 => x"20",
  2178 => x"20",
  2179 => x"20",
  2180 => x"00",
  2181 => x"3a",
  2182 => x"67",
  2183 => x"36",
  2184 => x"13",
  2185 => x"fc",
  2186 => x"00",
  2187 => x"10",
  2188 => x"00",
  2189 => x"7f",
  2190 => x"00",
  2191 => x"28",
  2192 => x"0c",
  2193 => x"a8",
  2194 => x"36",
  2195 => x"20",
  2196 => x"20",
  2197 => x"20",
  2198 => x"00",
  2199 => x"3a",
  2200 => x"67",
  2201 => x"24",
  2202 => x"13",
  2203 => x"fc",
  2204 => x"00",
  2205 => x"00",
  2206 => x"00",
  2207 => x"7f",
  2208 => x"00",
  2209 => x"28",
  2210 => x"0c",
  2211 => x"a8",
  2212 => x"46",
  2213 => x"41",
  2214 => x"54",
  2215 => x"33",
  2216 => x"00",
  2217 => x"52",
  2218 => x"66",
  2219 => x"ac",
  2220 => x"0c",
  2221 => x"a8",
  2222 => x"32",
  2223 => x"20",
  2224 => x"20",
  2225 => x"20",
  2226 => x"00",
  2227 => x"56",
  2228 => x"66",
  2229 => x"a2",
  2230 => x"13",
  2231 => x"fc",
  2232 => x"00",
  2233 => x"20",
  2234 => x"00",
  2235 => x"7f",
  2236 => x"00",
  2237 => x"28",
  2238 => x"20",
  2239 => x"28",
  2240 => x"00",
  2241 => x"0a",
  2242 => x"c0",
  2243 => x"bc",
  2244 => x"00",
  2245 => x"ff",
  2246 => x"ff",
  2247 => x"00",
  2248 => x"0c",
  2249 => x"80",
  2250 => x"00",
  2251 => x"00",
  2252 => x"02",
  2253 => x"00",
  2254 => x"66",
  2255 => x"88",
  2256 => x"22",
  2257 => x"39",
  2258 => x"00",
  2259 => x"7f",
  2260 => x"00",
  2261 => x"3e",
  2262 => x"30",
  2263 => x"28",
  2264 => x"00",
  2265 => x"0e",
  2266 => x"e0",
  2267 => x"58",
  2268 => x"d2",
  2269 => x"80",
  2270 => x"23",
  2271 => x"c1",
  2272 => x"00",
  2273 => x"7f",
  2274 => x"00",
  2275 => x"42",
  2276 => x"0c",
  2277 => x"39",
  2278 => x"00",
  2279 => x"20",
  2280 => x"00",
  2281 => x"7f",
  2282 => x"00",
  2283 => x"28",
  2284 => x"66",
  2285 => x"24",
  2286 => x"20",
  2287 => x"28",
  2288 => x"00",
  2289 => x"2c",
  2290 => x"e0",
  2291 => x"58",
  2292 => x"48",
  2293 => x"40",
  2294 => x"e0",
  2295 => x"58",
  2296 => x"23",
  2297 => x"c0",
  2298 => x"00",
  2299 => x"7f",
  2300 => x"00",
  2301 => x"2a",
  2302 => x"20",
  2303 => x"28",
  2304 => x"00",
  2305 => x"24",
  2306 => x"e0",
  2307 => x"58",
  2308 => x"48",
  2309 => x"40",
  2310 => x"e0",
  2311 => x"58",
  2312 => x"d2",
  2313 => x"80",
  2314 => x"53",
  2315 => x"28",
  2316 => x"00",
  2317 => x"10",
  2318 => x"66",
  2319 => x"f8",
  2320 => x"60",
  2321 => x"32",
  2322 => x"70",
  2323 => x"00",
  2324 => x"23",
  2325 => x"c0",
  2326 => x"00",
  2327 => x"7f",
  2328 => x"00",
  2329 => x"2a",
  2330 => x"30",
  2331 => x"28",
  2332 => x"00",
  2333 => x"16",
  2334 => x"e0",
  2335 => x"58",
  2336 => x"d2",
  2337 => x"80",
  2338 => x"53",
  2339 => x"28",
  2340 => x"00",
  2341 => x"10",
  2342 => x"66",
  2343 => x"f8",
  2344 => x"23",
  2345 => x"c1",
  2346 => x"00",
  2347 => x"7f",
  2348 => x"00",
  2349 => x"2e",
  2350 => x"20",
  2351 => x"01",
  2352 => x"10",
  2353 => x"28",
  2354 => x"00",
  2355 => x"12",
  2356 => x"e1",
  2357 => x"48",
  2358 => x"10",
  2359 => x"28",
  2360 => x"00",
  2361 => x"11",
  2362 => x"33",
  2363 => x"c0",
  2364 => x"00",
  2365 => x"7f",
  2366 => x"00",
  2367 => x"4e",
  2368 => x"e8",
  2369 => x"48",
  2370 => x"d2",
  2371 => x"80",
  2372 => x"70",
  2373 => x"00",
  2374 => x"10",
  2375 => x"28",
  2376 => x"00",
  2377 => x"0d",
  2378 => x"33",
  2379 => x"c0",
  2380 => x"00",
  2381 => x"7f",
  2382 => x"00",
  2383 => x"4a",
  2384 => x"92",
  2385 => x"80",
  2386 => x"92",
  2387 => x"80",
  2388 => x"23",
  2389 => x"c1",
  2390 => x"00",
  2391 => x"7f",
  2392 => x"00",
  2393 => x"46",
  2394 => x"33",
  2395 => x"fc",
  2396 => x"02",
  2397 => x"05",
  2398 => x"81",
  2399 => x"00",
  2400 => x"00",
  2401 => x"06",
  2402 => x"70",
  2403 => x"00",
  2404 => x"4e",
  2405 => x"75",
  2406 => x"20",
  2407 => x"39",
  2408 => x"00",
  2409 => x"7f",
  2410 => x"00",
  2411 => x"2a",
  2412 => x"23",
  2413 => x"c0",
  2414 => x"00",
  2415 => x"7f",
  2416 => x"00",
  2417 => x"32",
  2418 => x"66",
  2419 => x"28",
  2420 => x"42",
  2421 => x"b9",
  2422 => x"00",
  2423 => x"7f",
  2424 => x"00",
  2425 => x"32",
  2426 => x"30",
  2427 => x"39",
  2428 => x"00",
  2429 => x"7f",
  2430 => x"00",
  2431 => x"4e",
  2432 => x"e8",
  2433 => x"48",
  2434 => x"33",
  2435 => x"c0",
  2436 => x"00",
  2437 => x"7f",
  2438 => x"00",
  2439 => x"36",
  2440 => x"20",
  2441 => x"39",
  2442 => x"00",
  2443 => x"7f",
  2444 => x"00",
  2445 => x"2e",
  2446 => x"23",
  2447 => x"c0",
  2448 => x"00",
  2449 => x"7f",
  2450 => x"00",
  2451 => x"38",
  2452 => x"4e",
  2453 => x"75",
  2454 => x"20",
  2455 => x"39",
  2456 => x"00",
  2457 => x"7f",
  2458 => x"00",
  2459 => x"32",
  2460 => x"32",
  2461 => x"39",
  2462 => x"00",
  2463 => x"7f",
  2464 => x"00",
  2465 => x"4a",
  2466 => x"33",
  2467 => x"c1",
  2468 => x"00",
  2469 => x"7f",
  2470 => x"00",
  2471 => x"36",
  2472 => x"e2",
  2473 => x"49",
  2474 => x"65",
  2475 => x"04",
  2476 => x"e3",
  2477 => x"88",
  2478 => x"60",
  2479 => x"f8",
  2480 => x"d0",
  2481 => x"b9",
  2482 => x"00",
  2483 => x"7f",
  2484 => x"00",
  2485 => x"46",
  2486 => x"23",
  2487 => x"c0",
  2488 => x"00",
  2489 => x"7f",
  2490 => x"00",
  2491 => x"38",
  2492 => x"4e",
  2493 => x"75",
  2494 => x"48",
  2495 => x"e7",
  2496 => x"20",
  2497 => x"20",
  2498 => x"24",
  2499 => x"49",
  2500 => x"61",
  2501 => x"00",
  2502 => x"fa",
  2503 => x"10",
  2504 => x"66",
  2505 => x"7a",
  2506 => x"74",
  2507 => x"0f",
  2508 => x"4a",
  2509 => x"10",
  2510 => x"67",
  2511 => x"74",
  2512 => x"70",
  2513 => x"0a",
  2514 => x"12",
  2515 => x"32",
  2516 => x"00",
  2517 => x"00",
  2518 => x"b2",
  2519 => x"30",
  2520 => x"00",
  2521 => x"00",
  2522 => x"67",
  2523 => x"0a",
  2524 => x"d2",
  2525 => x"3c",
  2526 => x"00",
  2527 => x"20",
  2528 => x"b2",
  2529 => x"30",
  2530 => x"00",
  2531 => x"00",
  2532 => x"66",
  2533 => x"36",
  2534 => x"51",
  2535 => x"c8",
  2536 => x"ff",
  2537 => x"ea",
  2538 => x"70",
  2539 => x"00",
  2540 => x"10",
  2541 => x"28",
  2542 => x"00",
  2543 => x"0b",
  2544 => x"33",
  2545 => x"c0",
  2546 => x"00",
  2547 => x"7f",
  2548 => x"00",
  2549 => x"3c",
  2550 => x"0c",
  2551 => x"39",
  2552 => x"00",
  2553 => x"20",
  2554 => x"00",
  2555 => x"7f",
  2556 => x"00",
  2557 => x"28",
  2558 => x"66",
  2559 => x"08",
  2560 => x"30",
  2561 => x"28",
  2562 => x"00",
  2563 => x"14",
  2564 => x"e0",
  2565 => x"58",
  2566 => x"48",
  2567 => x"40",
  2568 => x"30",
  2569 => x"28",
  2570 => x"00",
  2571 => x"1a",
  2572 => x"e0",
  2573 => x"58",
  2574 => x"23",
  2575 => x"c0",
  2576 => x"00",
  2577 => x"7f",
  2578 => x"00",
  2579 => x"32",
  2580 => x"4c",
  2581 => x"df",
  2582 => x"04",
  2583 => x"04",
  2584 => x"70",
  2585 => x"ff",
  2586 => x"4e",
  2587 => x"75",
  2588 => x"41",
  2589 => x"e8",
  2590 => x"00",
  2591 => x"20",
  2592 => x"51",
  2593 => x"ca",
  2594 => x"ff",
  2595 => x"aa",
  2596 => x"20",
  2597 => x"39",
  2598 => x"00",
  2599 => x"7f",
  2600 => x"00",
  2601 => x"38",
  2602 => x"52",
  2603 => x"80",
  2604 => x"23",
  2605 => x"c0",
  2606 => x"00",
  2607 => x"7f",
  2608 => x"00",
  2609 => x"38",
  2610 => x"53",
  2611 => x"79",
  2612 => x"00",
  2613 => x"7f",
  2614 => x"00",
  2615 => x"36",
  2616 => x"66",
  2617 => x"8a",
  2618 => x"61",
  2619 => x"10",
  2620 => x"67",
  2621 => x"06",
  2622 => x"61",
  2623 => x"00",
  2624 => x"ff",
  2625 => x"56",
  2626 => x"60",
  2627 => x"80",
  2628 => x"4c",
  2629 => x"df",
  2630 => x"04",
  2631 => x"04",
  2632 => x"70",
  2633 => x"00",
  2634 => x"4e",
  2635 => x"75",
  2636 => x"0c",
  2637 => x"39",
  2638 => x"00",
  2639 => x"20",
  2640 => x"00",
  2641 => x"7f",
  2642 => x"00",
  2643 => x"28",
  2644 => x"67",
  2645 => x"3e",
  2646 => x"0c",
  2647 => x"39",
  2648 => x"00",
  2649 => x"0c",
  2650 => x"00",
  2651 => x"7f",
  2652 => x"00",
  2653 => x"28",
  2654 => x"67",
  2655 => x"78",
  2656 => x"20",
  2657 => x"39",
  2658 => x"00",
  2659 => x"7f",
  2660 => x"00",
  2661 => x"32",
  2662 => x"e0",
  2663 => x"88",
  2664 => x"d0",
  2665 => x"b9",
  2666 => x"00",
  2667 => x"7f",
  2668 => x"00",
  2669 => x"42",
  2670 => x"61",
  2671 => x"00",
  2672 => x"f9",
  2673 => x"66",
  2674 => x"66",
  2675 => x"60",
  2676 => x"10",
  2677 => x"39",
  2678 => x"00",
  2679 => x"7f",
  2680 => x"00",
  2681 => x"35",
  2682 => x"d0",
  2683 => x"40",
  2684 => x"30",
  2685 => x"30",
  2686 => x"00",
  2687 => x"00",
  2688 => x"e0",
  2689 => x"58",
  2690 => x"23",
  2691 => x"c0",
  2692 => x"00",
  2693 => x"7f",
  2694 => x"00",
  2695 => x"32",
  2696 => x"80",
  2697 => x"bc",
  2698 => x"ff",
  2699 => x"ff",
  2700 => x"00",
  2701 => x"0f",
  2702 => x"b0",
  2703 => x"7c",
  2704 => x"ff",
  2705 => x"ff",
  2706 => x"4e",
  2707 => x"75",
  2708 => x"20",
  2709 => x"39",
  2710 => x"00",
  2711 => x"7f",
  2712 => x"00",
  2713 => x"32",
  2714 => x"ee",
  2715 => x"88",
  2716 => x"d0",
  2717 => x"b9",
  2718 => x"00",
  2719 => x"7f",
  2720 => x"00",
  2721 => x"42",
  2722 => x"61",
  2723 => x"00",
  2724 => x"f9",
  2725 => x"32",
  2726 => x"66",
  2727 => x"2c",
  2728 => x"10",
  2729 => x"39",
  2730 => x"00",
  2731 => x"7f",
  2732 => x"00",
  2733 => x"35",
  2734 => x"c0",
  2735 => x"7c",
  2736 => x"00",
  2737 => x"7f",
  2738 => x"d0",
  2739 => x"40",
  2740 => x"d0",
  2741 => x"40",
  2742 => x"20",
  2743 => x"30",
  2744 => x"00",
  2745 => x"00",
  2746 => x"e0",
  2747 => x"58",
  2748 => x"48",
  2749 => x"40",
  2750 => x"e0",
  2751 => x"58",
  2752 => x"23",
  2753 => x"c0",
  2754 => x"00",
  2755 => x"7f",
  2756 => x"00",
  2757 => x"32",
  2758 => x"80",
  2759 => x"bc",
  2760 => x"f0",
  2761 => x"00",
  2762 => x"00",
  2763 => x"07",
  2764 => x"b0",
  2765 => x"bc",
  2766 => x"ff",
  2767 => x"ff",
  2768 => x"ff",
  2769 => x"ff",
  2770 => x"4e",
  2771 => x"75",
  2772 => x"70",
  2773 => x"00",
  2774 => x"4e",
  2775 => x"75",
  2776 => x"2f",
  2777 => x"02",
  2778 => x"20",
  2779 => x"39",
  2780 => x"00",
  2781 => x"7f",
  2782 => x"00",
  2783 => x"32",
  2784 => x"22",
  2785 => x"00",
  2786 => x"d0",
  2787 => x"80",
  2788 => x"d0",
  2789 => x"81",
  2790 => x"22",
  2791 => x"00",
  2792 => x"e0",
  2793 => x"88",
  2794 => x"e4",
  2795 => x"88",
  2796 => x"d0",
  2797 => x"b9",
  2798 => x"00",
  2799 => x"7f",
  2800 => x"00",
  2801 => x"42",
  2802 => x"24",
  2803 => x"00",
  2804 => x"61",
  2805 => x"00",
  2806 => x"f8",
  2807 => x"e0",
  2808 => x"66",
  2809 => x"52",
  2810 => x"20",
  2811 => x"01",
  2812 => x"e2",
  2813 => x"88",
  2814 => x"c0",
  2815 => x"7c",
  2816 => x"01",
  2817 => x"ff",
  2818 => x"b0",
  2819 => x"7c",
  2820 => x"01",
  2821 => x"ff",
  2822 => x"66",
  2823 => x"14",
  2824 => x"10",
  2825 => x"30",
  2826 => x"00",
  2827 => x"00",
  2828 => x"c1",
  2829 => x"42",
  2830 => x"52",
  2831 => x"80",
  2832 => x"61",
  2833 => x"00",
  2834 => x"f8",
  2835 => x"c4",
  2836 => x"66",
  2837 => x"36",
  2838 => x"e1",
  2839 => x"4a",
  2840 => x"14",
  2841 => x"10",
  2842 => x"60",
  2843 => x"0a",
  2844 => x"14",
  2845 => x"30",
  2846 => x"00",
  2847 => x"00",
  2848 => x"e1",
  2849 => x"4a",
  2850 => x"14",
  2851 => x"30",
  2852 => x"00",
  2853 => x"01",
  2854 => x"e1",
  2855 => x"5a",
  2856 => x"c2",
  2857 => x"7c",
  2858 => x"00",
  2859 => x"01",
  2860 => x"67",
  2861 => x"02",
  2862 => x"e8",
  2863 => x"4a",
  2864 => x"c4",
  2865 => x"bc",
  2866 => x"00",
  2867 => x"00",
  2868 => x"0f",
  2869 => x"ff",
  2870 => x"23",
  2871 => x"c2",
  2872 => x"00",
  2873 => x"7f",
  2874 => x"00",
  2875 => x"32",
  2876 => x"84",
  2877 => x"bc",
  2878 => x"ff",
  2879 => x"ff",
  2880 => x"f0",
  2881 => x"0f",
  2882 => x"20",
  2883 => x"02",
  2884 => x"24",
  2885 => x"1f",
  2886 => x"b0",
  2887 => x"7c",
  2888 => x"ff",
  2889 => x"ff",
  2890 => x"4e",
  2891 => x"75",
  2892 => x"24",
  2893 => x"1f",
  2894 => x"70",
  2895 => x"00",
  2896 => x"4e",
  2897 => x"75",
  2898 => x"41",
  2899 => x"f9",
  2900 => x"00",
  2901 => x"7f",
  2902 => x"00",
  2903 => x"04",
  2904 => x"20",
  2905 => x"bc",
  2906 => x"12",
  2907 => x"34",
  2908 => x"56",
  2909 => x"78",
  2910 => x"21",
  2911 => x"7c",
  2912 => x"fe",
  2913 => x"dc",
  2914 => x"ba",
  2915 => x"98",
  2916 => x"00",
  2917 => x"04",
  2918 => x"21",
  2919 => x"7c",
  2920 => x"aa",
  2921 => x"55",
  2922 => x"cc",
  2923 => x"22",
  2924 => x"00",
  2925 => x"02",
  2926 => x"11",
  2927 => x"7c",
  2928 => x"00",
  2929 => x"33",
  2930 => x"00",
  2931 => x"03",
  2932 => x"11",
  2933 => x"7c",
  2934 => x"00",
  2935 => x"fe",
  2936 => x"00",
  2937 => x"04",
  2938 => x"20",
  2939 => x"10",
  2940 => x"22",
  2941 => x"28",
  2942 => x"00",
  2943 => x"04",
  2944 => x"90",
  2945 => x"bc",
  2946 => x"12",
  2947 => x"34",
  2948 => x"aa",
  2949 => x"33",
  2950 => x"92",
  2951 => x"bc",
  2952 => x"fe",
  2953 => x"22",
  2954 => x"ba",
  2955 => x"98",
  2956 => x"80",
  2957 => x"81",
  2958 => x"4e",
  2959 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


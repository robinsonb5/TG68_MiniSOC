library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"41",
     9 => x"f9",
    10 => x"00",
    11 => x"10",
    12 => x"00",
    13 => x"00",
    14 => x"23",
    15 => x"c8",
    16 => x"80",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"70",
    21 => x"00",
    22 => x"2e",
    23 => x"3c",
    24 => x"00",
    25 => x"00",
    26 => x"01",
    27 => x"df",
    28 => x"2c",
    29 => x"3c",
    30 => x"00",
    31 => x"00",
    32 => x"02",
    33 => x"7f",
    34 => x"30",
    35 => x"c0",
    36 => x"52",
    37 => x"40",
    38 => x"51",
    39 => x"ce",
    40 => x"ff",
    41 => x"fa",
    42 => x"51",
    43 => x"cf",
    44 => x"ff",
    45 => x"f0",
    46 => x"41",
    47 => x"f9",
    48 => x"00",
    49 => x"10",
    50 => x"00",
    51 => x"00",
    52 => x"2e",
    53 => x"3c",
    54 => x"00",
    55 => x"00",
    56 => x"01",
    57 => x"df",
    58 => x"7c",
    59 => x"27",
    60 => x"4c",
    61 => x"d8",
    62 => x"1f",
    63 => x"1f",
    64 => x"51",
    65 => x"ce",
    66 => x"ff",
    67 => x"fa",
    68 => x"51",
    69 => x"cf",
    70 => x"ff",
    71 => x"f4",
    72 => x"60",
    73 => x"e4",
    74 => x"4f",
    75 => x"f9",
    76 => x"00",
    77 => x"7f",
    78 => x"00",
    79 => x"00",
    80 => x"70",
    81 => x"00",
    82 => x"30",
    83 => x"39",
    84 => x"81",
    85 => x"00",
    86 => x"00",
    87 => x"2a",
    88 => x"c0",
    89 => x"fc",
    90 => x"03",
    91 => x"e8",
    92 => x"80",
    93 => x"fc",
    94 => x"04",
    95 => x"80",
    96 => x"33",
    97 => x"c0",
    98 => x"81",
    99 => x"00",
   100 => x"00",
   101 => x"02",
   102 => x"46",
   103 => x"fc",
   104 => x"27",
   105 => x"00",
   106 => x"33",
   107 => x"fc",
   108 => x"f0",
   109 => x"00",
   110 => x"81",
   111 => x"00",
   112 => x"00",
   113 => x"06",
   114 => x"33",
   115 => x"fc",
   116 => x"00",
   117 => x"01",
   118 => x"81",
   119 => x"00",
   120 => x"00",
   121 => x"04",
   122 => x"41",
   123 => x"f9",
   124 => x"00",
   125 => x"7f",
   126 => x"00",
   127 => x"04",
   128 => x"20",
   129 => x"bc",
   130 => x"12",
   131 => x"34",
   132 => x"56",
   133 => x"78",
   134 => x"21",
   135 => x"7c",
   136 => x"fe",
   137 => x"dc",
   138 => x"ba",
   139 => x"98",
   140 => x"00",
   141 => x"04",
   142 => x"21",
   143 => x"7c",
   144 => x"aa",
   145 => x"55",
   146 => x"cc",
   147 => x"22",
   148 => x"00",
   149 => x"02",
   150 => x"11",
   151 => x"7c",
   152 => x"00",
   153 => x"33",
   154 => x"00",
   155 => x"03",
   156 => x"11",
   157 => x"7c",
   158 => x"00",
   159 => x"fe",
   160 => x"00",
   161 => x"04",
   162 => x"20",
   163 => x"10",
   164 => x"22",
   165 => x"28",
   166 => x"00",
   167 => x"04",
   168 => x"90",
   169 => x"bc",
   170 => x"12",
   171 => x"34",
   172 => x"aa",
   173 => x"33",
   174 => x"92",
   175 => x"bc",
   176 => x"fe",
   177 => x"22",
   178 => x"ba",
   179 => x"98",
   180 => x"41",
   181 => x"fa",
   182 => x"00",
   183 => x"74",
   184 => x"61",
   185 => x"00",
   186 => x"02",
   187 => x"d8",
   188 => x"33",
   189 => x"fc",
   190 => x"0f",
   191 => x"00",
   192 => x"81",
   193 => x"00",
   194 => x"00",
   195 => x"06",
   196 => x"2e",
   197 => x"3c",
   198 => x"00",
   199 => x"00",
   200 => x"07",
   201 => x"ff",
   202 => x"41",
   203 => x"f9",
   204 => x"80",
   205 => x"00",
   206 => x"08",
   207 => x"00",
   208 => x"10",
   209 => x"fc",
   210 => x"00",
   211 => x"20",
   212 => x"51",
   213 => x"cf",
   214 => x"ff",
   215 => x"fa",
   216 => x"23",
   217 => x"fc",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"7f",
   224 => x"00",
   225 => x"52",
   226 => x"41",
   227 => x"fa",
   228 => x"00",
   229 => x"46",
   230 => x"61",
   231 => x"00",
   232 => x"06",
   233 => x"ba",
   234 => x"61",
   235 => x"00",
   236 => x"0a",
   237 => x"ec",
   238 => x"4a",
   239 => x"80",
   240 => x"67",
   241 => x"0a",
   242 => x"41",
   243 => x"fa",
   244 => x"00",
   245 => x"6a",
   246 => x"61",
   247 => x"00",
   248 => x"06",
   249 => x"aa",
   250 => x"60",
   251 => x"fe",
   252 => x"41",
   253 => x"fa",
   254 => x"00",
   255 => x"49",
   256 => x"61",
   257 => x"00",
   258 => x"06",
   259 => x"a0",
   260 => x"61",
   261 => x"00",
   262 => x"02",
   263 => x"ac",
   264 => x"4b",
   265 => x"f9",
   266 => x"80",
   267 => x"00",
   268 => x"08",
   269 => x"00",
   270 => x"33",
   271 => x"fc",
   272 => x"00",
   273 => x"00",
   274 => x"00",
   275 => x"7f",
   276 => x"00",
   277 => x"0c",
   278 => x"30",
   279 => x"39",
   280 => x"81",
   281 => x"00",
   282 => x"00",
   283 => x"00",
   284 => x"08",
   285 => x"00",
   286 => x"00",
   287 => x"09",
   288 => x"67",
   289 => x"f4",
   290 => x"1a",
   291 => x"c0",
   292 => x"61",
   293 => x"00",
   294 => x"00",
   295 => x"80",
   296 => x"60",
   297 => x"ec",
   298 => x"43",
   299 => x"6f",
   300 => x"6e",
   301 => x"64",
   302 => x"75",
   303 => x"63",
   304 => x"74",
   305 => x"69",
   306 => x"6e",
   307 => x"67",
   308 => x"20",
   309 => x"73",
   310 => x"61",
   311 => x"6e",
   312 => x"69",
   313 => x"74",
   314 => x"79",
   315 => x"20",
   316 => x"63",
   317 => x"68",
   318 => x"65",
   319 => x"63",
   320 => x"6b",
   321 => x"2e",
   322 => x"2e",
   323 => x"2e",
   324 => x"0d",
   325 => x"0a",
   326 => x"00",
   327 => x"53",
   328 => x"61",
   329 => x"6e",
   330 => x"69",
   331 => x"74",
   332 => x"79",
   333 => x"20",
   334 => x"63",
   335 => x"68",
   336 => x"65",
   337 => x"63",
   338 => x"6b",
   339 => x"20",
   340 => x"70",
   341 => x"61",
   342 => x"73",
   343 => x"73",
   344 => x"65",
   345 => x"64",
   346 => x"2e",
   347 => x"0d",
   348 => x"0a",
   349 => x"00",
   350 => x"53",
   351 => x"61",
   352 => x"6e",
   353 => x"69",
   354 => x"74",
   355 => x"79",
   356 => x"20",
   357 => x"63",
   358 => x"68",
   359 => x"65",
   360 => x"63",
   361 => x"6b",
   362 => x"20",
   363 => x"66",
   364 => x"61",
   365 => x"69",
   366 => x"6c",
   367 => x"65",
   368 => x"64",
   369 => x"2e",
   370 => x"0d",
   371 => x"0a",
   372 => x"00",
   373 => x"00",
   374 => x"c0",
   375 => x"bc",
   376 => x"00",
   377 => x"00",
   378 => x"00",
   379 => x"df",
   380 => x"90",
   381 => x"3c",
   382 => x"00",
   383 => x"37",
   384 => x"6a",
   385 => x"04",
   386 => x"d0",
   387 => x"3c",
   388 => x"00",
   389 => x"27",
   390 => x"e9",
   391 => x"8e",
   392 => x"8c",
   393 => x"00",
   394 => x"20",
   395 => x"86",
   396 => x"4e",
   397 => x"75",
   398 => x"c0",
   399 => x"bc",
   400 => x"00",
   401 => x"00",
   402 => x"00",
   403 => x"df",
   404 => x"90",
   405 => x"3c",
   406 => x"00",
   407 => x"37",
   408 => x"6a",
   409 => x"04",
   410 => x"d0",
   411 => x"3c",
   412 => x"00",
   413 => x"27",
   414 => x"e9",
   415 => x"0f",
   416 => x"8e",
   417 => x"00",
   418 => x"10",
   419 => x"87",
   420 => x"4e",
   421 => x"75",
   422 => x"52",
   423 => x"79",
   424 => x"00",
   425 => x"7f",
   426 => x"00",
   427 => x"0c",
   428 => x"b0",
   429 => x"3c",
   430 => x"00",
   431 => x"53",
   432 => x"66",
   433 => x"2a",
   434 => x"33",
   435 => x"fc",
   436 => x"ff",
   437 => x"ff",
   438 => x"81",
   439 => x"00",
   440 => x"00",
   441 => x"06",
   442 => x"72",
   443 => x"00",
   444 => x"2e",
   445 => x"01",
   446 => x"2c",
   447 => x"01",
   448 => x"33",
   449 => x"c1",
   450 => x"00",
   451 => x"7f",
   452 => x"00",
   453 => x"0c",
   454 => x"23",
   455 => x"c1",
   456 => x"00",
   457 => x"7f",
   458 => x"00",
   459 => x"08",
   460 => x"23",
   461 => x"c1",
   462 => x"00",
   463 => x"7f",
   464 => x"00",
   465 => x"04",
   466 => x"23",
   467 => x"c1",
   468 => x"00",
   469 => x"7f",
   470 => x"00",
   471 => x"10",
   472 => x"60",
   473 => x"00",
   474 => x"01",
   475 => x"72",
   476 => x"2c",
   477 => x"39",
   478 => x"00",
   479 => x"7f",
   480 => x"00",
   481 => x"20",
   482 => x"2e",
   483 => x"39",
   484 => x"00",
   485 => x"7f",
   486 => x"00",
   487 => x"1c",
   488 => x"0c",
   489 => x"79",
   490 => x"00",
   491 => x"01",
   492 => x"00",
   493 => x"7f",
   494 => x"00",
   495 => x"0c",
   496 => x"66",
   497 => x"34",
   498 => x"33",
   499 => x"fc",
   500 => x"f0",
   501 => x"00",
   502 => x"81",
   503 => x"00",
   504 => x"00",
   505 => x"06",
   506 => x"41",
   507 => x"f9",
   508 => x"00",
   509 => x"7f",
   510 => x"00",
   511 => x"13",
   512 => x"61",
   513 => x"8c",
   514 => x"22",
   515 => x"39",
   516 => x"00",
   517 => x"7f",
   518 => x"00",
   519 => x"10",
   520 => x"b2",
   521 => x"bc",
   522 => x"00",
   523 => x"00",
   524 => x"00",
   525 => x"03",
   526 => x"6f",
   527 => x"08",
   528 => x"72",
   529 => x"0a",
   530 => x"92",
   531 => x"b9",
   532 => x"00",
   533 => x"7f",
   534 => x"00",
   535 => x"10",
   536 => x"52",
   537 => x"81",
   538 => x"e3",
   539 => x"89",
   540 => x"23",
   541 => x"c1",
   542 => x"00",
   543 => x"7f",
   544 => x"00",
   545 => x"14",
   546 => x"60",
   547 => x"00",
   548 => x"01",
   549 => x"28",
   550 => x"33",
   551 => x"f9",
   552 => x"00",
   553 => x"7f",
   554 => x"00",
   555 => x"12",
   556 => x"81",
   557 => x"00",
   558 => x"00",
   559 => x"06",
   560 => x"4a",
   561 => x"b9",
   562 => x"00",
   563 => x"7f",
   564 => x"00",
   565 => x"10",
   566 => x"67",
   567 => x"00",
   568 => x"01",
   569 => x"14",
   570 => x"0c",
   571 => x"b9",
   572 => x"00",
   573 => x"00",
   574 => x"00",
   575 => x"09",
   576 => x"00",
   577 => x"7f",
   578 => x"00",
   579 => x"10",
   580 => x"6e",
   581 => x"00",
   582 => x"00",
   583 => x"c0",
   584 => x"0c",
   585 => x"79",
   586 => x"00",
   587 => x"03",
   588 => x"00",
   589 => x"7f",
   590 => x"00",
   591 => x"0c",
   592 => x"6e",
   593 => x"16",
   594 => x"33",
   595 => x"fc",
   596 => x"0f",
   597 => x"00",
   598 => x"81",
   599 => x"00",
   600 => x"00",
   601 => x"06",
   602 => x"41",
   603 => x"f9",
   604 => x"00",
   605 => x"7f",
   606 => x"00",
   607 => x"07",
   608 => x"61",
   609 => x"00",
   610 => x"ff",
   611 => x"2c",
   612 => x"60",
   613 => x"00",
   614 => x"00",
   615 => x"e6",
   616 => x"22",
   617 => x"39",
   618 => x"00",
   619 => x"7f",
   620 => x"00",
   621 => x"14",
   622 => x"56",
   623 => x"41",
   624 => x"34",
   625 => x"39",
   626 => x"00",
   627 => x"7f",
   628 => x"00",
   629 => x"0c",
   630 => x"b4",
   631 => x"41",
   632 => x"6e",
   633 => x"20",
   634 => x"41",
   635 => x"f9",
   636 => x"00",
   637 => x"7f",
   638 => x"00",
   639 => x"08",
   640 => x"61",
   641 => x"00",
   642 => x"fe",
   643 => x"f4",
   644 => x"33",
   645 => x"f9",
   646 => x"00",
   647 => x"7f",
   648 => x"00",
   649 => x"0a",
   650 => x"81",
   651 => x"00",
   652 => x"00",
   653 => x"06",
   654 => x"33",
   655 => x"fc",
   656 => x"00",
   657 => x"01",
   658 => x"00",
   659 => x"7f",
   660 => x"00",
   661 => x"18",
   662 => x"60",
   663 => x"00",
   664 => x"00",
   665 => x"b4",
   666 => x"0c",
   667 => x"b9",
   668 => x"00",
   669 => x"00",
   670 => x"00",
   671 => x"03",
   672 => x"00",
   673 => x"7f",
   674 => x"00",
   675 => x"10",
   676 => x"6e",
   677 => x"60",
   678 => x"33",
   679 => x"fc",
   680 => x"00",
   681 => x"0f",
   682 => x"81",
   683 => x"00",
   684 => x"00",
   685 => x"06",
   686 => x"22",
   687 => x"39",
   688 => x"00",
   689 => x"7f",
   690 => x"00",
   691 => x"04",
   692 => x"e3",
   693 => x"89",
   694 => x"52",
   695 => x"81",
   696 => x"34",
   697 => x"39",
   698 => x"00",
   699 => x"7f",
   700 => x"00",
   701 => x"0c",
   702 => x"b4",
   703 => x"41",
   704 => x"6e",
   705 => x"2a",
   706 => x"20",
   707 => x"79",
   708 => x"00",
   709 => x"7f",
   710 => x"00",
   711 => x"08",
   712 => x"61",
   713 => x"00",
   714 => x"fe",
   715 => x"c4",
   716 => x"32",
   717 => x"39",
   718 => x"00",
   719 => x"7f",
   720 => x"00",
   721 => x"18",
   722 => x"53",
   723 => x"79",
   724 => x"00",
   725 => x"7f",
   726 => x"00",
   727 => x"18",
   728 => x"53",
   729 => x"41",
   730 => x"6a",
   731 => x"70",
   732 => x"52",
   733 => x"b9",
   734 => x"00",
   735 => x"7f",
   736 => x"00",
   737 => x"08",
   738 => x"33",
   739 => x"fc",
   740 => x"00",
   741 => x"01",
   742 => x"00",
   743 => x"7f",
   744 => x"00",
   745 => x"18",
   746 => x"60",
   747 => x"60",
   748 => x"30",
   749 => x"39",
   750 => x"00",
   751 => x"7f",
   752 => x"00",
   753 => x"18",
   754 => x"52",
   755 => x"40",
   756 => x"c0",
   757 => x"7c",
   758 => x"00",
   759 => x"01",
   760 => x"67",
   761 => x"52",
   762 => x"20",
   763 => x"79",
   764 => x"00",
   765 => x"7f",
   766 => x"00",
   767 => x"08",
   768 => x"e5",
   769 => x"88",
   770 => x"e1",
   771 => x"2f",
   772 => x"10",
   773 => x"87",
   774 => x"33",
   775 => x"fc",
   776 => x"f0",
   777 => x"f0",
   778 => x"81",
   779 => x"00",
   780 => x"00",
   781 => x"06",
   782 => x"0c",
   783 => x"b9",
   784 => x"00",
   785 => x"00",
   786 => x"00",
   787 => x"07",
   788 => x"00",
   789 => x"7f",
   790 => x"00",
   791 => x"10",
   792 => x"6d",
   793 => x"32",
   794 => x"33",
   795 => x"fc",
   796 => x"f0",
   797 => x"0f",
   798 => x"81",
   799 => x"00",
   800 => x"00",
   801 => x"06",
   802 => x"0c",
   803 => x"b9",
   804 => x"00",
   805 => x"00",
   806 => x"00",
   807 => x"09",
   808 => x"00",
   809 => x"7f",
   810 => x"00",
   811 => x"10",
   812 => x"6e",
   813 => x"1e",
   814 => x"33",
   815 => x"fc",
   816 => x"ff",
   817 => x"f0",
   818 => x"81",
   819 => x"00",
   820 => x"00",
   821 => x"06",
   822 => x"41",
   823 => x"fa",
   824 => x"00",
   825 => x"22",
   826 => x"61",
   827 => x"56",
   828 => x"2e",
   829 => x"b9",
   830 => x"00",
   831 => x"7f",
   832 => x"00",
   833 => x"08",
   834 => x"08",
   835 => x"b9",
   836 => x"00",
   837 => x"00",
   838 => x"81",
   839 => x"00",
   840 => x"00",
   841 => x"04",
   842 => x"4e",
   843 => x"75",
   844 => x"23",
   845 => x"c6",
   846 => x"00",
   847 => x"7f",
   848 => x"00",
   849 => x"20",
   850 => x"23",
   851 => x"c7",
   852 => x"00",
   853 => x"7f",
   854 => x"00",
   855 => x"1c",
   856 => x"4e",
   857 => x"75",
   858 => x"46",
   859 => x"69",
   860 => x"72",
   861 => x"6d",
   862 => x"77",
   863 => x"61",
   864 => x"72",
   865 => x"65",
   866 => x"20",
   867 => x"72",
   868 => x"65",
   869 => x"63",
   870 => x"65",
   871 => x"69",
   872 => x"76",
   873 => x"65",
   874 => x"64",
   875 => x"20",
   876 => x"2d",
   877 => x"20",
   878 => x"6c",
   879 => x"61",
   880 => x"75",
   881 => x"6e",
   882 => x"63",
   883 => x"68",
   884 => x"69",
   885 => x"6e",
   886 => x"67",
   887 => x"0d",
   888 => x"0a",
   889 => x"00",
   890 => x"48",
   891 => x"40",
   892 => x"30",
   893 => x"39",
   894 => x"81",
   895 => x"00",
   896 => x"00",
   897 => x"00",
   898 => x"08",
   899 => x"00",
   900 => x"00",
   901 => x"08",
   902 => x"67",
   903 => x"f4",
   904 => x"48",
   905 => x"40",
   906 => x"33",
   907 => x"c0",
   908 => x"81",
   909 => x"00",
   910 => x"00",
   911 => x"00",
   912 => x"4e",
   913 => x"75",
   914 => x"2f",
   915 => x"00",
   916 => x"70",
   917 => x"00",
   918 => x"30",
   919 => x"39",
   920 => x"81",
   921 => x"00",
   922 => x"00",
   923 => x"00",
   924 => x"08",
   925 => x"00",
   926 => x"00",
   927 => x"08",
   928 => x"67",
   929 => x"f4",
   930 => x"10",
   931 => x"18",
   932 => x"67",
   933 => x"08",
   934 => x"33",
   935 => x"c0",
   936 => x"81",
   937 => x"00",
   938 => x"00",
   939 => x"00",
   940 => x"60",
   941 => x"e8",
   942 => x"20",
   943 => x"1f",
   944 => x"4e",
   945 => x"75",
   946 => x"33",
   947 => x"fc",
   948 => x"00",
   949 => x"01",
   950 => x"81",
   951 => x"00",
   952 => x"00",
   953 => x"06",
   954 => x"41",
   955 => x"fa",
   956 => x"01",
   957 => x"fa",
   958 => x"61",
   959 => x"00",
   960 => x"03",
   961 => x"e2",
   962 => x"61",
   963 => x"00",
   964 => x"02",
   965 => x"60",
   966 => x"66",
   967 => x"5c",
   968 => x"33",
   969 => x"fc",
   970 => x"00",
   971 => x"02",
   972 => x"81",
   973 => x"00",
   974 => x"00",
   975 => x"06",
   976 => x"33",
   977 => x"fc",
   978 => x"00",
   979 => x"40",
   980 => x"00",
   981 => x"7f",
   982 => x"00",
   983 => x"26",
   984 => x"61",
   985 => x"00",
   986 => x"04",
   987 => x"8a",
   988 => x"67",
   989 => x"0c",
   990 => x"42",
   991 => x"79",
   992 => x"00",
   993 => x"7f",
   994 => x"00",
   995 => x"26",
   996 => x"61",
   997 => x"00",
   998 => x"04",
   999 => x"7e",
  1000 => x"66",
  1001 => x"28",
  1002 => x"33",
  1003 => x"fc",
  1004 => x"00",
  1005 => x"03",
  1006 => x"81",
  1007 => x"00",
  1008 => x"00",
  1009 => x"06",
  1010 => x"61",
  1011 => x"00",
  1012 => x"05",
  1013 => x"f8",
  1014 => x"43",
  1015 => x"fa",
  1016 => x"00",
  1017 => x"57",
  1018 => x"61",
  1019 => x"00",
  1020 => x"06",
  1021 => x"48",
  1022 => x"67",
  1023 => x"12",
  1024 => x"41",
  1025 => x"fa",
  1026 => x"00",
  1027 => x"47",
  1028 => x"61",
  1029 => x"00",
  1030 => x"03",
  1031 => x"9c",
  1032 => x"30",
  1033 => x"7c",
  1034 => x"20",
  1035 => x"00",
  1036 => x"61",
  1037 => x"00",
  1038 => x"04",
  1039 => x"02",
  1040 => x"4e",
  1041 => x"75",
  1042 => x"33",
  1043 => x"fc",
  1044 => x"f0",
  1045 => x"03",
  1046 => x"81",
  1047 => x"00",
  1048 => x"00",
  1049 => x"06",
  1050 => x"41",
  1051 => x"fa",
  1052 => x"00",
  1053 => x"29",
  1054 => x"61",
  1055 => x"00",
  1056 => x"03",
  1057 => x"82",
  1058 => x"4e",
  1059 => x"75",
  1060 => x"33",
  1061 => x"fc",
  1062 => x"f0",
  1063 => x"02",
  1064 => x"81",
  1065 => x"00",
  1066 => x"00",
  1067 => x"06",
  1068 => x"41",
  1069 => x"fa",
  1070 => x"00",
  1071 => x"08",
  1072 => x"61",
  1073 => x"00",
  1074 => x"03",
  1075 => x"70",
  1076 => x"4e",
  1077 => x"75",
  1078 => x"53",
  1079 => x"44",
  1080 => x"20",
  1081 => x"69",
  1082 => x"6e",
  1083 => x"69",
  1084 => x"74",
  1085 => x"20",
  1086 => x"66",
  1087 => x"61",
  1088 => x"69",
  1089 => x"6c",
  1090 => x"65",
  1091 => x"64",
  1092 => x"00",
  1093 => x"6e",
  1094 => x"6f",
  1095 => x"74",
  1096 => x"20",
  1097 => x"66",
  1098 => x"6f",
  1099 => x"75",
  1100 => x"6e",
  1101 => x"64",
  1102 => x"20",
  1103 => x"42",
  1104 => x"4f",
  1105 => x"4f",
  1106 => x"54",
  1107 => x"20",
  1108 => x"20",
  1109 => x"20",
  1110 => x"20",
  1111 => x"53",
  1112 => x"52",
  1113 => x"45",
  1114 => x"00",
  1115 => x"00",
  1116 => x"33",
  1117 => x"fc",
  1118 => x"01",
  1119 => x"00",
  1120 => x"81",
  1121 => x"00",
  1122 => x"00",
  1123 => x"06",
  1124 => x"41",
  1125 => x"f9",
  1126 => x"00",
  1127 => x"7f",
  1128 => x"00",
  1129 => x"56",
  1130 => x"61",
  1131 => x"00",
  1132 => x"00",
  1133 => x"c4",
  1134 => x"66",
  1135 => x"68",
  1136 => x"33",
  1137 => x"fc",
  1138 => x"01",
  1139 => x"01",
  1140 => x"81",
  1141 => x"00",
  1142 => x"00",
  1143 => x"06",
  1144 => x"32",
  1145 => x"3c",
  1146 => x"4e",
  1147 => x"20",
  1148 => x"53",
  1149 => x"41",
  1150 => x"67",
  1151 => x"44",
  1152 => x"33",
  1153 => x"fc",
  1154 => x"01",
  1155 => x"02",
  1156 => x"81",
  1157 => x"00",
  1158 => x"00",
  1159 => x"06",
  1160 => x"33",
  1161 => x"7c",
  1162 => x"00",
  1163 => x"ff",
  1164 => x"00",
  1165 => x"24",
  1166 => x"30",
  1167 => x"29",
  1168 => x"00",
  1169 => x"24",
  1170 => x"b0",
  1171 => x"3c",
  1172 => x"00",
  1173 => x"fe",
  1174 => x"66",
  1175 => x"e4",
  1176 => x"30",
  1177 => x"29",
  1178 => x"01",
  1179 => x"00",
  1180 => x"32",
  1181 => x"3c",
  1182 => x"00",
  1183 => x"7f",
  1184 => x"20",
  1185 => x"29",
  1186 => x"01",
  1187 => x"00",
  1188 => x"20",
  1189 => x"c0",
  1190 => x"51",
  1191 => x"c9",
  1192 => x"ff",
  1193 => x"f8",
  1194 => x"30",
  1195 => x"29",
  1196 => x"00",
  1197 => x"24",
  1198 => x"33",
  1199 => x"7c",
  1200 => x"00",
  1201 => x"00",
  1202 => x"00",
  1203 => x"22",
  1204 => x"33",
  1205 => x"fc",
  1206 => x"01",
  1207 => x"03",
  1208 => x"81",
  1209 => x"00",
  1210 => x"00",
  1211 => x"06",
  1212 => x"41",
  1213 => x"e8",
  1214 => x"fe",
  1215 => x"00",
  1216 => x"70",
  1217 => x"00",
  1218 => x"4e",
  1219 => x"75",
  1220 => x"33",
  1221 => x"fc",
  1222 => x"f1",
  1223 => x"02",
  1224 => x"81",
  1225 => x"00",
  1226 => x"00",
  1227 => x"06",
  1228 => x"41",
  1229 => x"fa",
  1230 => x"01",
  1231 => x"38",
  1232 => x"61",
  1233 => x"00",
  1234 => x"02",
  1235 => x"d0",
  1236 => x"70",
  1237 => x"fe",
  1238 => x"4e",
  1239 => x"75",
  1240 => x"33",
  1241 => x"fc",
  1242 => x"f1",
  1243 => x"03",
  1244 => x"81",
  1245 => x"00",
  1246 => x"00",
  1247 => x"06",
  1248 => x"41",
  1249 => x"fa",
  1250 => x"01",
  1251 => x"0c",
  1252 => x"61",
  1253 => x"00",
  1254 => x"02",
  1255 => x"bc",
  1256 => x"70",
  1257 => x"ff",
  1258 => x"4e",
  1259 => x"75",
  1260 => x"22",
  1261 => x"3c",
  1262 => x"00",
  1263 => x"95",
  1264 => x"00",
  1265 => x"40",
  1266 => x"70",
  1267 => x"00",
  1268 => x"60",
  1269 => x"40",
  1270 => x"22",
  1271 => x"3c",
  1272 => x"00",
  1273 => x"ff",
  1274 => x"00",
  1275 => x"41",
  1276 => x"70",
  1277 => x"00",
  1278 => x"60",
  1279 => x"36",
  1280 => x"22",
  1281 => x"3c",
  1282 => x"00",
  1283 => x"87",
  1284 => x"00",
  1285 => x"48",
  1286 => x"20",
  1287 => x"3c",
  1288 => x"00",
  1289 => x"00",
  1290 => x"01",
  1291 => x"aa",
  1292 => x"60",
  1293 => x"28",
  1294 => x"22",
  1295 => x"3c",
  1296 => x"00",
  1297 => x"87",
  1298 => x"00",
  1299 => x"69",
  1300 => x"20",
  1301 => x"3c",
  1302 => x"40",
  1303 => x"00",
  1304 => x"00",
  1305 => x"00",
  1306 => x"60",
  1307 => x"1a",
  1308 => x"22",
  1309 => x"3c",
  1310 => x"00",
  1311 => x"ff",
  1312 => x"00",
  1313 => x"77",
  1314 => x"70",
  1315 => x"00",
  1316 => x"60",
  1317 => x"10",
  1318 => x"22",
  1319 => x"3c",
  1320 => x"00",
  1321 => x"ff",
  1322 => x"00",
  1323 => x"7a",
  1324 => x"70",
  1325 => x"00",
  1326 => x"60",
  1327 => x"06",
  1328 => x"22",
  1329 => x"3c",
  1330 => x"00",
  1331 => x"ff",
  1332 => x"00",
  1333 => x"51",
  1334 => x"43",
  1335 => x"f9",
  1336 => x"81",
  1337 => x"00",
  1338 => x"00",
  1339 => x"00",
  1340 => x"33",
  1341 => x"7c",
  1342 => x"00",
  1343 => x"ff",
  1344 => x"00",
  1345 => x"24",
  1346 => x"3f",
  1347 => x"69",
  1348 => x"00",
  1349 => x"24",
  1350 => x"ff",
  1351 => x"fe",
  1352 => x"33",
  1353 => x"7c",
  1354 => x"00",
  1355 => x"01",
  1356 => x"00",
  1357 => x"22",
  1358 => x"33",
  1359 => x"7c",
  1360 => x"00",
  1361 => x"ff",
  1362 => x"00",
  1363 => x"24",
  1364 => x"33",
  1365 => x"41",
  1366 => x"00",
  1367 => x"24",
  1368 => x"48",
  1369 => x"41",
  1370 => x"4a",
  1371 => x"79",
  1372 => x"00",
  1373 => x"7f",
  1374 => x"00",
  1375 => x"24",
  1376 => x"67",
  1377 => x"16",
  1378 => x"e1",
  1379 => x"98",
  1380 => x"33",
  1381 => x"40",
  1382 => x"00",
  1383 => x"24",
  1384 => x"e1",
  1385 => x"98",
  1386 => x"33",
  1387 => x"40",
  1388 => x"00",
  1389 => x"24",
  1390 => x"e1",
  1391 => x"98",
  1392 => x"33",
  1393 => x"40",
  1394 => x"00",
  1395 => x"24",
  1396 => x"e1",
  1397 => x"98",
  1398 => x"60",
  1399 => x"18",
  1400 => x"d0",
  1401 => x"80",
  1402 => x"48",
  1403 => x"40",
  1404 => x"33",
  1405 => x"40",
  1406 => x"00",
  1407 => x"24",
  1408 => x"48",
  1409 => x"40",
  1410 => x"e1",
  1411 => x"58",
  1412 => x"33",
  1413 => x"40",
  1414 => x"00",
  1415 => x"24",
  1416 => x"e1",
  1417 => x"58",
  1418 => x"33",
  1419 => x"40",
  1420 => x"00",
  1421 => x"24",
  1422 => x"70",
  1423 => x"00",
  1424 => x"33",
  1425 => x"40",
  1426 => x"00",
  1427 => x"24",
  1428 => x"33",
  1429 => x"41",
  1430 => x"00",
  1431 => x"24",
  1432 => x"22",
  1433 => x"3c",
  1434 => x"00",
  1435 => x"00",
  1436 => x"01",
  1437 => x"90",
  1438 => x"53",
  1439 => x"81",
  1440 => x"67",
  1441 => x"10",
  1442 => x"33",
  1443 => x"7c",
  1444 => x"00",
  1445 => x"ff",
  1446 => x"00",
  1447 => x"24",
  1448 => x"30",
  1449 => x"29",
  1450 => x"00",
  1451 => x"24",
  1452 => x"b0",
  1453 => x"3c",
  1454 => x"00",
  1455 => x"ff",
  1456 => x"67",
  1457 => x"ec",
  1458 => x"80",
  1459 => x"00",
  1460 => x"4e",
  1461 => x"75",
  1462 => x"53",
  1463 => x"74",
  1464 => x"61",
  1465 => x"72",
  1466 => x"74",
  1467 => x"20",
  1468 => x"49",
  1469 => x"6e",
  1470 => x"69",
  1471 => x"74",
  1472 => x"0d",
  1473 => x"0a",
  1474 => x"00",
  1475 => x"49",
  1476 => x"6e",
  1477 => x"69",
  1478 => x"74",
  1479 => x"20",
  1480 => x"64",
  1481 => x"6f",
  1482 => x"6e",
  1483 => x"65",
  1484 => x"0d",
  1485 => x"0a",
  1486 => x"00",
  1487 => x"49",
  1488 => x"6e",
  1489 => x"69",
  1490 => x"74",
  1491 => x"20",
  1492 => x"66",
  1493 => x"61",
  1494 => x"69",
  1495 => x"6c",
  1496 => x"75",
  1497 => x"72",
  1498 => x"65",
  1499 => x"0d",
  1500 => x"0a",
  1501 => x"00",
  1502 => x"52",
  1503 => x"65",
  1504 => x"73",
  1505 => x"65",
  1506 => x"74",
  1507 => x"20",
  1508 => x"66",
  1509 => x"61",
  1510 => x"69",
  1511 => x"6c",
  1512 => x"75",
  1513 => x"72",
  1514 => x"65",
  1515 => x"0d",
  1516 => x"0a",
  1517 => x"00",
  1518 => x"43",
  1519 => x"6f",
  1520 => x"6d",
  1521 => x"6d",
  1522 => x"61",
  1523 => x"6e",
  1524 => x"64",
  1525 => x"20",
  1526 => x"54",
  1527 => x"69",
  1528 => x"6d",
  1529 => x"65",
  1530 => x"6f",
  1531 => x"75",
  1532 => x"74",
  1533 => x"5f",
  1534 => x"45",
  1535 => x"72",
  1536 => x"72",
  1537 => x"6f",
  1538 => x"72",
  1539 => x"0d",
  1540 => x"0a",
  1541 => x"00",
  1542 => x"54",
  1543 => x"69",
  1544 => x"6d",
  1545 => x"65",
  1546 => x"6f",
  1547 => x"75",
  1548 => x"74",
  1549 => x"5f",
  1550 => x"45",
  1551 => x"72",
  1552 => x"72",
  1553 => x"6f",
  1554 => x"72",
  1555 => x"0d",
  1556 => x"0a",
  1557 => x"00",
  1558 => x"53",
  1559 => x"44",
  1560 => x"48",
  1561 => x"43",
  1562 => x"20",
  1563 => x"66",
  1564 => x"6f",
  1565 => x"75",
  1566 => x"6e",
  1567 => x"64",
  1568 => x"20",
  1569 => x"0d",
  1570 => x"0a",
  1571 => x"00",
  1572 => x"33",
  1573 => x"fc",
  1574 => x"ff",
  1575 => x"ff",
  1576 => x"00",
  1577 => x"7f",
  1578 => x"00",
  1579 => x"24",
  1580 => x"43",
  1581 => x"f9",
  1582 => x"81",
  1583 => x"00",
  1584 => x"00",
  1585 => x"00",
  1586 => x"33",
  1587 => x"7c",
  1588 => x"00",
  1589 => x"00",
  1590 => x"00",
  1591 => x"22",
  1592 => x"33",
  1593 => x"7c",
  1594 => x"00",
  1595 => x"96",
  1596 => x"00",
  1597 => x"1e",
  1598 => x"32",
  1599 => x"3c",
  1600 => x"00",
  1601 => x"c8",
  1602 => x"43",
  1603 => x"e9",
  1604 => x"00",
  1605 => x"20",
  1606 => x"33",
  1607 => x"7c",
  1608 => x"00",
  1609 => x"ff",
  1610 => x"00",
  1611 => x"24",
  1612 => x"51",
  1613 => x"c9",
  1614 => x"ff",
  1615 => x"f8",
  1616 => x"34",
  1617 => x"3c",
  1618 => x"00",
  1619 => x"32",
  1620 => x"61",
  1621 => x"00",
  1622 => x"fe",
  1623 => x"96",
  1624 => x"3f",
  1625 => x"69",
  1626 => x"00",
  1627 => x"24",
  1628 => x"ff",
  1629 => x"fe",
  1630 => x"33",
  1631 => x"7c",
  1632 => x"00",
  1633 => x"00",
  1634 => x"00",
  1635 => x"22",
  1636 => x"b0",
  1637 => x"3c",
  1638 => x"00",
  1639 => x"01",
  1640 => x"67",
  1641 => x"12",
  1642 => x"51",
  1643 => x"ca",
  1644 => x"ff",
  1645 => x"e8",
  1646 => x"48",
  1647 => x"7a",
  1648 => x"ff",
  1649 => x"6e",
  1650 => x"61",
  1651 => x"00",
  1652 => x"01",
  1653 => x"22",
  1654 => x"58",
  1655 => x"8f",
  1656 => x"70",
  1657 => x"ff",
  1658 => x"4e",
  1659 => x"75",
  1660 => x"22",
  1661 => x"3c",
  1662 => x"00",
  1663 => x"00",
  1664 => x"20",
  1665 => x"00",
  1666 => x"33",
  1667 => x"7c",
  1668 => x"00",
  1669 => x"ff",
  1670 => x"00",
  1671 => x"24",
  1672 => x"53",
  1673 => x"81",
  1674 => x"66",
  1675 => x"f6",
  1676 => x"61",
  1677 => x"00",
  1678 => x"fe",
  1679 => x"72",
  1680 => x"b0",
  1681 => x"3c",
  1682 => x"00",
  1683 => x"01",
  1684 => x"66",
  1685 => x"00",
  1686 => x"00",
  1687 => x"9e",
  1688 => x"33",
  1689 => x"7c",
  1690 => x"00",
  1691 => x"ff",
  1692 => x"00",
  1693 => x"24",
  1694 => x"33",
  1695 => x"7c",
  1696 => x"00",
  1697 => x"ff",
  1698 => x"00",
  1699 => x"24",
  1700 => x"33",
  1701 => x"7c",
  1702 => x"00",
  1703 => x"ff",
  1704 => x"00",
  1705 => x"24",
  1706 => x"30",
  1707 => x"29",
  1708 => x"00",
  1709 => x"24",
  1710 => x"0c",
  1711 => x"00",
  1712 => x"00",
  1713 => x"01",
  1714 => x"66",
  1715 => x"00",
  1716 => x"00",
  1717 => x"80",
  1718 => x"33",
  1719 => x"7c",
  1720 => x"00",
  1721 => x"ff",
  1722 => x"00",
  1723 => x"24",
  1724 => x"30",
  1725 => x"29",
  1726 => x"00",
  1727 => x"24",
  1728 => x"0c",
  1729 => x"00",
  1730 => x"00",
  1731 => x"aa",
  1732 => x"66",
  1733 => x"6e",
  1734 => x"3f",
  1735 => x"69",
  1736 => x"00",
  1737 => x"24",
  1738 => x"ff",
  1739 => x"fe",
  1740 => x"33",
  1741 => x"7c",
  1742 => x"00",
  1743 => x"00",
  1744 => x"00",
  1745 => x"22",
  1746 => x"48",
  1747 => x"7a",
  1748 => x"ff",
  1749 => x"42",
  1750 => x"61",
  1751 => x"00",
  1752 => x"00",
  1753 => x"be",
  1754 => x"58",
  1755 => x"8f",
  1756 => x"34",
  1757 => x"3c",
  1758 => x"00",
  1759 => x"32",
  1760 => x"53",
  1761 => x"42",
  1762 => x"67",
  1763 => x"50",
  1764 => x"32",
  1765 => x"3c",
  1766 => x"07",
  1767 => x"d0",
  1768 => x"33",
  1769 => x"7c",
  1770 => x"00",
  1771 => x"ff",
  1772 => x"00",
  1773 => x"24",
  1774 => x"51",
  1775 => x"c9",
  1776 => x"ff",
  1777 => x"f8",
  1778 => x"61",
  1779 => x"00",
  1780 => x"fe",
  1781 => x"28",
  1782 => x"b0",
  1783 => x"3c",
  1784 => x"00",
  1785 => x"01",
  1786 => x"66",
  1787 => x"e4",
  1788 => x"61",
  1789 => x"00",
  1790 => x"fe",
  1791 => x"10",
  1792 => x"66",
  1793 => x"de",
  1794 => x"61",
  1795 => x"00",
  1796 => x"fe",
  1797 => x"22",
  1798 => x"66",
  1799 => x"d8",
  1800 => x"33",
  1801 => x"7c",
  1802 => x"00",
  1803 => x"ff",
  1804 => x"00",
  1805 => x"24",
  1806 => x"30",
  1807 => x"29",
  1808 => x"00",
  1809 => x"24",
  1810 => x"c0",
  1811 => x"3c",
  1812 => x"00",
  1813 => x"40",
  1814 => x"66",
  1815 => x"08",
  1816 => x"33",
  1817 => x"fc",
  1818 => x"00",
  1819 => x"00",
  1820 => x"00",
  1821 => x"7f",
  1822 => x"00",
  1823 => x"24",
  1824 => x"33",
  1825 => x"7c",
  1826 => x"00",
  1827 => x"ff",
  1828 => x"00",
  1829 => x"24",
  1830 => x"33",
  1831 => x"7c",
  1832 => x"00",
  1833 => x"ff",
  1834 => x"00",
  1835 => x"24",
  1836 => x"33",
  1837 => x"7c",
  1838 => x"00",
  1839 => x"ff",
  1840 => x"00",
  1841 => x"24",
  1842 => x"60",
  1843 => x"3c",
  1844 => x"33",
  1845 => x"fc",
  1846 => x"00",
  1847 => x"00",
  1848 => x"00",
  1849 => x"7f",
  1850 => x"00",
  1851 => x"24",
  1852 => x"34",
  1853 => x"3c",
  1854 => x"00",
  1855 => x"0a",
  1856 => x"32",
  1857 => x"3c",
  1858 => x"07",
  1859 => x"d0",
  1860 => x"33",
  1861 => x"7c",
  1862 => x"00",
  1863 => x"ff",
  1864 => x"00",
  1865 => x"24",
  1866 => x"51",
  1867 => x"c9",
  1868 => x"ff",
  1869 => x"f8",
  1870 => x"61",
  1871 => x"00",
  1872 => x"fd",
  1873 => x"a6",
  1874 => x"67",
  1875 => x"1c",
  1876 => x"3f",
  1877 => x"69",
  1878 => x"00",
  1879 => x"24",
  1880 => x"ff",
  1881 => x"fe",
  1882 => x"33",
  1883 => x"7c",
  1884 => x"00",
  1885 => x"00",
  1886 => x"00",
  1887 => x"22",
  1888 => x"51",
  1889 => x"ca",
  1890 => x"ff",
  1891 => x"de",
  1892 => x"48",
  1893 => x"7a",
  1894 => x"fe",
  1895 => x"69",
  1896 => x"61",
  1897 => x"2c",
  1898 => x"58",
  1899 => x"8f",
  1900 => x"70",
  1901 => x"ff",
  1902 => x"4e",
  1903 => x"75",
  1904 => x"3f",
  1905 => x"69",
  1906 => x"00",
  1907 => x"24",
  1908 => x"ff",
  1909 => x"fe",
  1910 => x"33",
  1911 => x"7c",
  1912 => x"00",
  1913 => x"00",
  1914 => x"00",
  1915 => x"22",
  1916 => x"33",
  1917 => x"69",
  1918 => x"00",
  1919 => x"2c",
  1920 => x"00",
  1921 => x"1e",
  1922 => x"48",
  1923 => x"7a",
  1924 => x"fe",
  1925 => x"3f",
  1926 => x"61",
  1927 => x"0e",
  1928 => x"58",
  1929 => x"8f",
  1930 => x"33",
  1931 => x"fc",
  1932 => x"ff",
  1933 => x"ff",
  1934 => x"81",
  1935 => x"00",
  1936 => x"00",
  1937 => x"06",
  1938 => x"70",
  1939 => x"00",
  1940 => x"4e",
  1941 => x"75",
  1942 => x"2f",
  1943 => x"08",
  1944 => x"20",
  1945 => x"6f",
  1946 => x"00",
  1947 => x"08",
  1948 => x"61",
  1949 => x"04",
  1950 => x"20",
  1951 => x"5f",
  1952 => x"4e",
  1953 => x"75",
  1954 => x"48",
  1955 => x"e7",
  1956 => x"00",
  1957 => x"c0",
  1958 => x"22",
  1959 => x"39",
  1960 => x"00",
  1961 => x"7f",
  1962 => x"00",
  1963 => x"52",
  1964 => x"43",
  1965 => x"f9",
  1966 => x"80",
  1967 => x"00",
  1968 => x"08",
  1969 => x"00",
  1970 => x"10",
  1971 => x"18",
  1972 => x"67",
  1973 => x"08",
  1974 => x"13",
  1975 => x"80",
  1976 => x"10",
  1977 => x"00",
  1978 => x"52",
  1979 => x"41",
  1980 => x"60",
  1981 => x"f4",
  1982 => x"06",
  1983 => x"b9",
  1984 => x"00",
  1985 => x"00",
  1986 => x"00",
  1987 => x"4c",
  1988 => x"00",
  1989 => x"7f",
  1990 => x"00",
  1991 => x"52",
  1992 => x"4c",
  1993 => x"df",
  1994 => x"03",
  1995 => x"00",
  1996 => x"4e",
  1997 => x"75",
  1998 => x"4a",
  1999 => x"79",
  2000 => x"00",
  2001 => x"7f",
  2002 => x"00",
  2003 => x"24",
  2004 => x"67",
  2005 => x"1e",
  2006 => x"41",
  2007 => x"fa",
  2008 => x"00",
  2009 => x"08",
  2010 => x"48",
  2011 => x"7a",
  2012 => x"00",
  2013 => x"34",
  2014 => x"60",
  2015 => x"c2",
  2016 => x"53",
  2017 => x"44",
  2018 => x"48",
  2019 => x"43",
  2020 => x"20",
  2021 => x"66",
  2022 => x"6c",
  2023 => x"61",
  2024 => x"67",
  2025 => x"20",
  2026 => x"73",
  2027 => x"74",
  2028 => x"69",
  2029 => x"6c",
  2030 => x"6c",
  2031 => x"20",
  2032 => x"73",
  2033 => x"65",
  2034 => x"74",
  2035 => x"00",
  2036 => x"41",
  2037 => x"fa",
  2038 => x"00",
  2039 => x"08",
  2040 => x"48",
  2041 => x"7a",
  2042 => x"00",
  2043 => x"16",
  2044 => x"60",
  2045 => x"a4",
  2046 => x"53",
  2047 => x"44",
  2048 => x"48",
  2049 => x"43",
  2050 => x"20",
  2051 => x"66",
  2052 => x"6c",
  2053 => x"61",
  2054 => x"67",
  2055 => x"20",
  2056 => x"63",
  2057 => x"6c",
  2058 => x"65",
  2059 => x"61",
  2060 => x"72",
  2061 => x"65",
  2062 => x"64",
  2063 => x"00",
  2064 => x"61",
  2065 => x"00",
  2066 => x"02",
  2067 => x"0a",
  2068 => x"61",
  2069 => x"00",
  2070 => x"fc",
  2071 => x"46",
  2072 => x"66",
  2073 => x"46",
  2074 => x"2e",
  2075 => x"3c",
  2076 => x"00",
  2077 => x"00",
  2078 => x"01",
  2079 => x"ff",
  2080 => x"41",
  2081 => x"f9",
  2082 => x"00",
  2083 => x"7f",
  2084 => x"00",
  2085 => x"56",
  2086 => x"43",
  2087 => x"f9",
  2088 => x"80",
  2089 => x"00",
  2090 => x"08",
  2091 => x"00",
  2092 => x"10",
  2093 => x"18",
  2094 => x"12",
  2095 => x"c0",
  2096 => x"48",
  2097 => x"e7",
  2098 => x"01",
  2099 => x"c0",
  2100 => x"61",
  2101 => x"00",
  2102 => x"f9",
  2103 => x"70",
  2104 => x"4c",
  2105 => x"df",
  2106 => x"03",
  2107 => x"80",
  2108 => x"51",
  2109 => x"cf",
  2110 => x"ff",
  2111 => x"ee",
  2112 => x"20",
  2113 => x"39",
  2114 => x"00",
  2115 => x"7f",
  2116 => x"00",
  2117 => x"38",
  2118 => x"52",
  2119 => x"80",
  2120 => x"23",
  2121 => x"c0",
  2122 => x"00",
  2123 => x"7f",
  2124 => x"00",
  2125 => x"38",
  2126 => x"53",
  2127 => x"79",
  2128 => x"00",
  2129 => x"7f",
  2130 => x"00",
  2131 => x"36",
  2132 => x"66",
  2133 => x"be",
  2134 => x"61",
  2135 => x"00",
  2136 => x"02",
  2137 => x"7a",
  2138 => x"66",
  2139 => x"b4",
  2140 => x"20",
  2141 => x"08",
  2142 => x"4e",
  2143 => x"75",
  2144 => x"70",
  2145 => x"00",
  2146 => x"4e",
  2147 => x"75",
  2148 => x"33",
  2149 => x"fc",
  2150 => x"02",
  2151 => x"01",
  2152 => x"81",
  2153 => x"00",
  2154 => x"00",
  2155 => x"06",
  2156 => x"70",
  2157 => x"00",
  2158 => x"23",
  2159 => x"c0",
  2160 => x"00",
  2161 => x"7f",
  2162 => x"00",
  2163 => x"3e",
  2164 => x"33",
  2165 => x"fc",
  2166 => x"02",
  2167 => x"11",
  2168 => x"81",
  2169 => x"00",
  2170 => x"00",
  2171 => x"06",
  2172 => x"61",
  2173 => x"00",
  2174 => x"fb",
  2175 => x"de",
  2176 => x"66",
  2177 => x"5c",
  2178 => x"33",
  2179 => x"fc",
  2180 => x"02",
  2181 => x"02",
  2182 => x"81",
  2183 => x"00",
  2184 => x"00",
  2185 => x"06",
  2186 => x"0c",
  2187 => x"28",
  2188 => x"00",
  2189 => x"55",
  2190 => x"01",
  2191 => x"fe",
  2192 => x"66",
  2193 => x"4c",
  2194 => x"0c",
  2195 => x"28",
  2196 => x"00",
  2197 => x"aa",
  2198 => x"01",
  2199 => x"ff",
  2200 => x"66",
  2201 => x"44",
  2202 => x"30",
  2203 => x"39",
  2204 => x"00",
  2205 => x"7f",
  2206 => x"00",
  2207 => x"26",
  2208 => x"c0",
  2209 => x"7c",
  2210 => x"00",
  2211 => x"70",
  2212 => x"b0",
  2213 => x"7c",
  2214 => x"00",
  2215 => x"40",
  2216 => x"64",
  2217 => x"40",
  2218 => x"43",
  2219 => x"e8",
  2220 => x"01",
  2221 => x"be",
  2222 => x"d2",
  2223 => x"c0",
  2224 => x"33",
  2225 => x"fc",
  2226 => x"02",
  2227 => x"03",
  2228 => x"81",
  2229 => x"00",
  2230 => x"00",
  2231 => x"06",
  2232 => x"20",
  2233 => x"29",
  2234 => x"00",
  2235 => x"08",
  2236 => x"e0",
  2237 => x"58",
  2238 => x"48",
  2239 => x"40",
  2240 => x"e0",
  2241 => x"58",
  2242 => x"23",
  2243 => x"c0",
  2244 => x"00",
  2245 => x"7f",
  2246 => x"00",
  2247 => x"3e",
  2248 => x"61",
  2249 => x"00",
  2250 => x"fb",
  2251 => x"92",
  2252 => x"66",
  2253 => x"10",
  2254 => x"0c",
  2255 => x"28",
  2256 => x"00",
  2257 => x"55",
  2258 => x"01",
  2259 => x"fe",
  2260 => x"66",
  2261 => x"08",
  2262 => x"0c",
  2263 => x"28",
  2264 => x"00",
  2265 => x"aa",
  2266 => x"01",
  2267 => x"ff",
  2268 => x"67",
  2269 => x"0c",
  2270 => x"33",
  2271 => x"fc",
  2272 => x"f2",
  2273 => x"01",
  2274 => x"81",
  2275 => x"00",
  2276 => x"00",
  2277 => x"06",
  2278 => x"70",
  2279 => x"ff",
  2280 => x"4e",
  2281 => x"75",
  2282 => x"33",
  2283 => x"fc",
  2284 => x"02",
  2285 => x"04",
  2286 => x"81",
  2287 => x"00",
  2288 => x"00",
  2289 => x"06",
  2290 => x"0c",
  2291 => x"a8",
  2292 => x"46",
  2293 => x"41",
  2294 => x"54",
  2295 => x"31",
  2296 => x"00",
  2297 => x"36",
  2298 => x"66",
  2299 => x"24",
  2300 => x"13",
  2301 => x"fc",
  2302 => x"00",
  2303 => x"0c",
  2304 => x"00",
  2305 => x"7f",
  2306 => x"00",
  2307 => x"28",
  2308 => x"0c",
  2309 => x"a8",
  2310 => x"32",
  2311 => x"20",
  2312 => x"20",
  2313 => x"20",
  2314 => x"00",
  2315 => x"3a",
  2316 => x"67",
  2317 => x"36",
  2318 => x"13",
  2319 => x"fc",
  2320 => x"00",
  2321 => x"10",
  2322 => x"00",
  2323 => x"7f",
  2324 => x"00",
  2325 => x"28",
  2326 => x"0c",
  2327 => x"a8",
  2328 => x"36",
  2329 => x"20",
  2330 => x"20",
  2331 => x"20",
  2332 => x"00",
  2333 => x"3a",
  2334 => x"67",
  2335 => x"24",
  2336 => x"13",
  2337 => x"fc",
  2338 => x"00",
  2339 => x"00",
  2340 => x"00",
  2341 => x"7f",
  2342 => x"00",
  2343 => x"28",
  2344 => x"0c",
  2345 => x"a8",
  2346 => x"46",
  2347 => x"41",
  2348 => x"54",
  2349 => x"33",
  2350 => x"00",
  2351 => x"52",
  2352 => x"66",
  2353 => x"ac",
  2354 => x"0c",
  2355 => x"a8",
  2356 => x"32",
  2357 => x"20",
  2358 => x"20",
  2359 => x"20",
  2360 => x"00",
  2361 => x"56",
  2362 => x"66",
  2363 => x"a2",
  2364 => x"13",
  2365 => x"fc",
  2366 => x"00",
  2367 => x"20",
  2368 => x"00",
  2369 => x"7f",
  2370 => x"00",
  2371 => x"28",
  2372 => x"20",
  2373 => x"28",
  2374 => x"00",
  2375 => x"0a",
  2376 => x"c0",
  2377 => x"bc",
  2378 => x"00",
  2379 => x"ff",
  2380 => x"ff",
  2381 => x"00",
  2382 => x"0c",
  2383 => x"80",
  2384 => x"00",
  2385 => x"00",
  2386 => x"02",
  2387 => x"00",
  2388 => x"66",
  2389 => x"88",
  2390 => x"22",
  2391 => x"39",
  2392 => x"00",
  2393 => x"7f",
  2394 => x"00",
  2395 => x"3e",
  2396 => x"30",
  2397 => x"28",
  2398 => x"00",
  2399 => x"0e",
  2400 => x"e0",
  2401 => x"58",
  2402 => x"d2",
  2403 => x"80",
  2404 => x"23",
  2405 => x"c1",
  2406 => x"00",
  2407 => x"7f",
  2408 => x"00",
  2409 => x"42",
  2410 => x"0c",
  2411 => x"39",
  2412 => x"00",
  2413 => x"20",
  2414 => x"00",
  2415 => x"7f",
  2416 => x"00",
  2417 => x"28",
  2418 => x"66",
  2419 => x"24",
  2420 => x"20",
  2421 => x"28",
  2422 => x"00",
  2423 => x"2c",
  2424 => x"e0",
  2425 => x"58",
  2426 => x"48",
  2427 => x"40",
  2428 => x"e0",
  2429 => x"58",
  2430 => x"23",
  2431 => x"c0",
  2432 => x"00",
  2433 => x"7f",
  2434 => x"00",
  2435 => x"2a",
  2436 => x"20",
  2437 => x"28",
  2438 => x"00",
  2439 => x"24",
  2440 => x"e0",
  2441 => x"58",
  2442 => x"48",
  2443 => x"40",
  2444 => x"e0",
  2445 => x"58",
  2446 => x"d2",
  2447 => x"80",
  2448 => x"53",
  2449 => x"28",
  2450 => x"00",
  2451 => x"10",
  2452 => x"66",
  2453 => x"f8",
  2454 => x"60",
  2455 => x"32",
  2456 => x"70",
  2457 => x"00",
  2458 => x"23",
  2459 => x"c0",
  2460 => x"00",
  2461 => x"7f",
  2462 => x"00",
  2463 => x"2a",
  2464 => x"30",
  2465 => x"28",
  2466 => x"00",
  2467 => x"16",
  2468 => x"e0",
  2469 => x"58",
  2470 => x"d2",
  2471 => x"80",
  2472 => x"53",
  2473 => x"28",
  2474 => x"00",
  2475 => x"10",
  2476 => x"66",
  2477 => x"f8",
  2478 => x"23",
  2479 => x"c1",
  2480 => x"00",
  2481 => x"7f",
  2482 => x"00",
  2483 => x"2e",
  2484 => x"20",
  2485 => x"01",
  2486 => x"10",
  2487 => x"28",
  2488 => x"00",
  2489 => x"12",
  2490 => x"e1",
  2491 => x"48",
  2492 => x"10",
  2493 => x"28",
  2494 => x"00",
  2495 => x"11",
  2496 => x"33",
  2497 => x"c0",
  2498 => x"00",
  2499 => x"7f",
  2500 => x"00",
  2501 => x"4e",
  2502 => x"e8",
  2503 => x"48",
  2504 => x"d2",
  2505 => x"80",
  2506 => x"70",
  2507 => x"00",
  2508 => x"10",
  2509 => x"28",
  2510 => x"00",
  2511 => x"0d",
  2512 => x"33",
  2513 => x"c0",
  2514 => x"00",
  2515 => x"7f",
  2516 => x"00",
  2517 => x"4a",
  2518 => x"92",
  2519 => x"80",
  2520 => x"92",
  2521 => x"80",
  2522 => x"23",
  2523 => x"c1",
  2524 => x"00",
  2525 => x"7f",
  2526 => x"00",
  2527 => x"46",
  2528 => x"33",
  2529 => x"fc",
  2530 => x"02",
  2531 => x"05",
  2532 => x"81",
  2533 => x"00",
  2534 => x"00",
  2535 => x"06",
  2536 => x"70",
  2537 => x"00",
  2538 => x"4e",
  2539 => x"75",
  2540 => x"20",
  2541 => x"39",
  2542 => x"00",
  2543 => x"7f",
  2544 => x"00",
  2545 => x"2a",
  2546 => x"23",
  2547 => x"c0",
  2548 => x"00",
  2549 => x"7f",
  2550 => x"00",
  2551 => x"32",
  2552 => x"66",
  2553 => x"28",
  2554 => x"42",
  2555 => x"b9",
  2556 => x"00",
  2557 => x"7f",
  2558 => x"00",
  2559 => x"32",
  2560 => x"30",
  2561 => x"39",
  2562 => x"00",
  2563 => x"7f",
  2564 => x"00",
  2565 => x"4e",
  2566 => x"e8",
  2567 => x"48",
  2568 => x"33",
  2569 => x"c0",
  2570 => x"00",
  2571 => x"7f",
  2572 => x"00",
  2573 => x"36",
  2574 => x"20",
  2575 => x"39",
  2576 => x"00",
  2577 => x"7f",
  2578 => x"00",
  2579 => x"2e",
  2580 => x"23",
  2581 => x"c0",
  2582 => x"00",
  2583 => x"7f",
  2584 => x"00",
  2585 => x"38",
  2586 => x"4e",
  2587 => x"75",
  2588 => x"20",
  2589 => x"39",
  2590 => x"00",
  2591 => x"7f",
  2592 => x"00",
  2593 => x"32",
  2594 => x"32",
  2595 => x"39",
  2596 => x"00",
  2597 => x"7f",
  2598 => x"00",
  2599 => x"4a",
  2600 => x"33",
  2601 => x"c1",
  2602 => x"00",
  2603 => x"7f",
  2604 => x"00",
  2605 => x"36",
  2606 => x"e2",
  2607 => x"49",
  2608 => x"65",
  2609 => x"04",
  2610 => x"e3",
  2611 => x"88",
  2612 => x"60",
  2613 => x"f8",
  2614 => x"d0",
  2615 => x"b9",
  2616 => x"00",
  2617 => x"7f",
  2618 => x"00",
  2619 => x"46",
  2620 => x"23",
  2621 => x"c0",
  2622 => x"00",
  2623 => x"7f",
  2624 => x"00",
  2625 => x"38",
  2626 => x"4e",
  2627 => x"75",
  2628 => x"48",
  2629 => x"e7",
  2630 => x"20",
  2631 => x"20",
  2632 => x"24",
  2633 => x"49",
  2634 => x"61",
  2635 => x"00",
  2636 => x"fa",
  2637 => x"10",
  2638 => x"66",
  2639 => x"7a",
  2640 => x"74",
  2641 => x"0f",
  2642 => x"4a",
  2643 => x"10",
  2644 => x"67",
  2645 => x"74",
  2646 => x"70",
  2647 => x"0a",
  2648 => x"12",
  2649 => x"32",
  2650 => x"00",
  2651 => x"00",
  2652 => x"b2",
  2653 => x"30",
  2654 => x"00",
  2655 => x"00",
  2656 => x"67",
  2657 => x"0a",
  2658 => x"d2",
  2659 => x"3c",
  2660 => x"00",
  2661 => x"20",
  2662 => x"b2",
  2663 => x"30",
  2664 => x"00",
  2665 => x"00",
  2666 => x"66",
  2667 => x"36",
  2668 => x"51",
  2669 => x"c8",
  2670 => x"ff",
  2671 => x"ea",
  2672 => x"70",
  2673 => x"00",
  2674 => x"10",
  2675 => x"28",
  2676 => x"00",
  2677 => x"0b",
  2678 => x"33",
  2679 => x"c0",
  2680 => x"00",
  2681 => x"7f",
  2682 => x"00",
  2683 => x"3c",
  2684 => x"0c",
  2685 => x"39",
  2686 => x"00",
  2687 => x"20",
  2688 => x"00",
  2689 => x"7f",
  2690 => x"00",
  2691 => x"28",
  2692 => x"66",
  2693 => x"08",
  2694 => x"30",
  2695 => x"28",
  2696 => x"00",
  2697 => x"14",
  2698 => x"e0",
  2699 => x"58",
  2700 => x"48",
  2701 => x"40",
  2702 => x"30",
  2703 => x"28",
  2704 => x"00",
  2705 => x"1a",
  2706 => x"e0",
  2707 => x"58",
  2708 => x"23",
  2709 => x"c0",
  2710 => x"00",
  2711 => x"7f",
  2712 => x"00",
  2713 => x"32",
  2714 => x"4c",
  2715 => x"df",
  2716 => x"04",
  2717 => x"04",
  2718 => x"70",
  2719 => x"ff",
  2720 => x"4e",
  2721 => x"75",
  2722 => x"41",
  2723 => x"e8",
  2724 => x"00",
  2725 => x"20",
  2726 => x"51",
  2727 => x"ca",
  2728 => x"ff",
  2729 => x"aa",
  2730 => x"20",
  2731 => x"39",
  2732 => x"00",
  2733 => x"7f",
  2734 => x"00",
  2735 => x"38",
  2736 => x"52",
  2737 => x"80",
  2738 => x"23",
  2739 => x"c0",
  2740 => x"00",
  2741 => x"7f",
  2742 => x"00",
  2743 => x"38",
  2744 => x"53",
  2745 => x"79",
  2746 => x"00",
  2747 => x"7f",
  2748 => x"00",
  2749 => x"36",
  2750 => x"66",
  2751 => x"8a",
  2752 => x"61",
  2753 => x"10",
  2754 => x"67",
  2755 => x"06",
  2756 => x"61",
  2757 => x"00",
  2758 => x"ff",
  2759 => x"56",
  2760 => x"60",
  2761 => x"80",
  2762 => x"4c",
  2763 => x"df",
  2764 => x"04",
  2765 => x"04",
  2766 => x"70",
  2767 => x"00",
  2768 => x"4e",
  2769 => x"75",
  2770 => x"0c",
  2771 => x"39",
  2772 => x"00",
  2773 => x"20",
  2774 => x"00",
  2775 => x"7f",
  2776 => x"00",
  2777 => x"28",
  2778 => x"67",
  2779 => x"3e",
  2780 => x"0c",
  2781 => x"39",
  2782 => x"00",
  2783 => x"0c",
  2784 => x"00",
  2785 => x"7f",
  2786 => x"00",
  2787 => x"28",
  2788 => x"67",
  2789 => x"78",
  2790 => x"20",
  2791 => x"39",
  2792 => x"00",
  2793 => x"7f",
  2794 => x"00",
  2795 => x"32",
  2796 => x"e0",
  2797 => x"88",
  2798 => x"d0",
  2799 => x"b9",
  2800 => x"00",
  2801 => x"7f",
  2802 => x"00",
  2803 => x"42",
  2804 => x"61",
  2805 => x"00",
  2806 => x"f9",
  2807 => x"66",
  2808 => x"66",
  2809 => x"60",
  2810 => x"10",
  2811 => x"39",
  2812 => x"00",
  2813 => x"7f",
  2814 => x"00",
  2815 => x"35",
  2816 => x"d0",
  2817 => x"40",
  2818 => x"30",
  2819 => x"30",
  2820 => x"00",
  2821 => x"00",
  2822 => x"e0",
  2823 => x"58",
  2824 => x"23",
  2825 => x"c0",
  2826 => x"00",
  2827 => x"7f",
  2828 => x"00",
  2829 => x"32",
  2830 => x"80",
  2831 => x"bc",
  2832 => x"ff",
  2833 => x"ff",
  2834 => x"00",
  2835 => x"0f",
  2836 => x"b0",
  2837 => x"7c",
  2838 => x"ff",
  2839 => x"ff",
  2840 => x"4e",
  2841 => x"75",
  2842 => x"20",
  2843 => x"39",
  2844 => x"00",
  2845 => x"7f",
  2846 => x"00",
  2847 => x"32",
  2848 => x"ee",
  2849 => x"88",
  2850 => x"d0",
  2851 => x"b9",
  2852 => x"00",
  2853 => x"7f",
  2854 => x"00",
  2855 => x"42",
  2856 => x"61",
  2857 => x"00",
  2858 => x"f9",
  2859 => x"32",
  2860 => x"66",
  2861 => x"2c",
  2862 => x"10",
  2863 => x"39",
  2864 => x"00",
  2865 => x"7f",
  2866 => x"00",
  2867 => x"35",
  2868 => x"c0",
  2869 => x"7c",
  2870 => x"00",
  2871 => x"7f",
  2872 => x"d0",
  2873 => x"40",
  2874 => x"d0",
  2875 => x"40",
  2876 => x"20",
  2877 => x"30",
  2878 => x"00",
  2879 => x"00",
  2880 => x"e0",
  2881 => x"58",
  2882 => x"48",
  2883 => x"40",
  2884 => x"e0",
  2885 => x"58",
  2886 => x"23",
  2887 => x"c0",
  2888 => x"00",
  2889 => x"7f",
  2890 => x"00",
  2891 => x"32",
  2892 => x"80",
  2893 => x"bc",
  2894 => x"f0",
  2895 => x"00",
  2896 => x"00",
  2897 => x"07",
  2898 => x"b0",
  2899 => x"bc",
  2900 => x"ff",
  2901 => x"ff",
  2902 => x"ff",
  2903 => x"ff",
  2904 => x"4e",
  2905 => x"75",
  2906 => x"70",
  2907 => x"00",
  2908 => x"4e",
  2909 => x"75",
  2910 => x"2f",
  2911 => x"02",
  2912 => x"20",
  2913 => x"39",
  2914 => x"00",
  2915 => x"7f",
  2916 => x"00",
  2917 => x"32",
  2918 => x"22",
  2919 => x"00",
  2920 => x"d0",
  2921 => x"80",
  2922 => x"d0",
  2923 => x"81",
  2924 => x"22",
  2925 => x"00",
  2926 => x"e0",
  2927 => x"88",
  2928 => x"e4",
  2929 => x"88",
  2930 => x"d0",
  2931 => x"b9",
  2932 => x"00",
  2933 => x"7f",
  2934 => x"00",
  2935 => x"42",
  2936 => x"24",
  2937 => x"00",
  2938 => x"61",
  2939 => x"00",
  2940 => x"f8",
  2941 => x"e0",
  2942 => x"66",
  2943 => x"52",
  2944 => x"20",
  2945 => x"01",
  2946 => x"e2",
  2947 => x"88",
  2948 => x"c0",
  2949 => x"7c",
  2950 => x"01",
  2951 => x"ff",
  2952 => x"b0",
  2953 => x"7c",
  2954 => x"01",
  2955 => x"ff",
  2956 => x"66",
  2957 => x"14",
  2958 => x"10",
  2959 => x"30",
  2960 => x"00",
  2961 => x"00",
  2962 => x"c1",
  2963 => x"42",
  2964 => x"52",
  2965 => x"80",
  2966 => x"61",
  2967 => x"00",
  2968 => x"f8",
  2969 => x"c4",
  2970 => x"66",
  2971 => x"36",
  2972 => x"e1",
  2973 => x"4a",
  2974 => x"14",
  2975 => x"10",
  2976 => x"60",
  2977 => x"0a",
  2978 => x"14",
  2979 => x"30",
  2980 => x"00",
  2981 => x"00",
  2982 => x"e1",
  2983 => x"4a",
  2984 => x"14",
  2985 => x"30",
  2986 => x"00",
  2987 => x"01",
  2988 => x"e1",
  2989 => x"5a",
  2990 => x"c2",
  2991 => x"7c",
  2992 => x"00",
  2993 => x"01",
  2994 => x"67",
  2995 => x"02",
  2996 => x"e8",
  2997 => x"4a",
  2998 => x"c4",
  2999 => x"bc",
  3000 => x"00",
  3001 => x"00",
  3002 => x"0f",
  3003 => x"ff",
  3004 => x"23",
  3005 => x"c2",
  3006 => x"00",
  3007 => x"7f",
  3008 => x"00",
  3009 => x"32",
  3010 => x"84",
  3011 => x"bc",
  3012 => x"ff",
  3013 => x"ff",
  3014 => x"f0",
  3015 => x"0f",
  3016 => x"20",
  3017 => x"02",
  3018 => x"24",
  3019 => x"1f",
  3020 => x"b0",
  3021 => x"7c",
  3022 => x"ff",
  3023 => x"ff",
  3024 => x"4e",
  3025 => x"75",
  3026 => x"24",
  3027 => x"1f",
  3028 => x"70",
  3029 => x"00",
  3030 => x"4e",
  3031 => x"75",
  3032 => x"41",
  3033 => x"f9",
  3034 => x"00",
  3035 => x"7f",
  3036 => x"00",
  3037 => x"04",
  3038 => x"20",
  3039 => x"bc",
  3040 => x"12",
  3041 => x"34",
  3042 => x"56",
  3043 => x"78",
  3044 => x"21",
  3045 => x"7c",
  3046 => x"fe",
  3047 => x"dc",
  3048 => x"ba",
  3049 => x"98",
  3050 => x"00",
  3051 => x"04",
  3052 => x"21",
  3053 => x"7c",
  3054 => x"aa",
  3055 => x"55",
  3056 => x"cc",
  3057 => x"22",
  3058 => x"00",
  3059 => x"02",
  3060 => x"11",
  3061 => x"7c",
  3062 => x"00",
  3063 => x"33",
  3064 => x"00",
  3065 => x"03",
  3066 => x"11",
  3067 => x"7c",
  3068 => x"00",
  3069 => x"fe",
  3070 => x"00",
  3071 => x"04",
  3072 => x"20",
  3073 => x"10",
  3074 => x"22",
  3075 => x"28",
  3076 => x"00",
  3077 => x"04",
  3078 => x"90",
  3079 => x"bc",
  3080 => x"12",
  3081 => x"34",
  3082 => x"aa",
  3083 => x"33",
  3084 => x"92",
  3085 => x"bc",
  3086 => x"fe",
  3087 => x"22",
  3088 => x"ba",
  3089 => x"98",
  3090 => x"80",
  3091 => x"81",
  3092 => x"4e",
  3093 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


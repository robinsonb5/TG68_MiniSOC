library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SanityCheck_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end SanityCheck_ROM;

architecture arch of SanityCheck_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"00",
     2 => x"0f",
     3 => x"fe",
     4 => x"00",
     5 => x"00",
     6 => x"01",
     7 => x"00",
     8 => x"00",
     9 => x"00",
    10 => x"00",
    11 => x"00",
    12 => x"00",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"00",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"00",
    21 => x"00",
    22 => x"00",
    23 => x"00",
    24 => x"00",
    25 => x"00",
    26 => x"00",
    27 => x"00",
    28 => x"00",
    29 => x"00",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"00",
    34 => x"00",
    35 => x"00",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"00",
    40 => x"00",
    41 => x"00",
    42 => x"00",
    43 => x"00",
    44 => x"00",
    45 => x"00",
    46 => x"00",
    47 => x"00",
    48 => x"00",
    49 => x"00",
    50 => x"00",
    51 => x"00",
    52 => x"00",
    53 => x"00",
    54 => x"00",
    55 => x"00",
    56 => x"00",
    57 => x"00",
    58 => x"00",
    59 => x"00",
    60 => x"00",
    61 => x"00",
    62 => x"00",
    63 => x"00",
    64 => x"00",
    65 => x"00",
    66 => x"00",
    67 => x"00",
    68 => x"00",
    69 => x"00",
    70 => x"00",
    71 => x"00",
    72 => x"00",
    73 => x"00",
    74 => x"00",
    75 => x"00",
    76 => x"00",
    77 => x"00",
    78 => x"00",
    79 => x"00",
    80 => x"00",
    81 => x"00",
    82 => x"00",
    83 => x"00",
    84 => x"00",
    85 => x"00",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"00",
    93 => x"00",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"00",
   127 => x"00",
   128 => x"00",
   129 => x"00",
   130 => x"00",
   131 => x"00",
   132 => x"00",
   133 => x"00",
   134 => x"00",
   135 => x"00",
   136 => x"00",
   137 => x"00",
   138 => x"00",
   139 => x"00",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"00",
   144 => x"00",
   145 => x"00",
   146 => x"00",
   147 => x"00",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"00",
   153 => x"00",
   154 => x"00",
   155 => x"00",
   156 => x"00",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"00",
   161 => x"00",
   162 => x"00",
   163 => x"00",
   164 => x"00",
   165 => x"00",
   166 => x"00",
   167 => x"00",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"00",
   172 => x"00",
   173 => x"00",
   174 => x"00",
   175 => x"00",
   176 => x"00",
   177 => x"00",
   178 => x"00",
   179 => x"00",
   180 => x"00",
   181 => x"00",
   182 => x"00",
   183 => x"00",
   184 => x"00",
   185 => x"00",
   186 => x"00",
   187 => x"00",
   188 => x"00",
   189 => x"00",
   190 => x"00",
   191 => x"00",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"00",
   196 => x"00",
   197 => x"00",
   198 => x"00",
   199 => x"00",
   200 => x"00",
   201 => x"00",
   202 => x"00",
   203 => x"00",
   204 => x"00",
   205 => x"00",
   206 => x"00",
   207 => x"00",
   208 => x"00",
   209 => x"00",
   210 => x"00",
   211 => x"00",
   212 => x"00",
   213 => x"00",
   214 => x"00",
   215 => x"00",
   216 => x"00",
   217 => x"00",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"00",
   224 => x"00",
   225 => x"00",
   226 => x"00",
   227 => x"00",
   228 => x"00",
   229 => x"00",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"00",
   234 => x"00",
   235 => x"00",
   236 => x"00",
   237 => x"00",
   238 => x"00",
   239 => x"00",
   240 => x"00",
   241 => x"00",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"00",
   248 => x"00",
   249 => x"00",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"00",
   256 => x"4f",
   257 => x"f9",
   258 => x"00",
   259 => x"00",
   260 => x"0f",
   261 => x"fe",
   262 => x"41",
   263 => x"f9",
   264 => x"00",
   265 => x"00",
   266 => x"0b",
   267 => x"6c",
   268 => x"20",
   269 => x"3c",
   270 => x"00",
   271 => x"00",
   272 => x"0b",
   273 => x"6c",
   274 => x"b1",
   275 => x"c0",
   276 => x"6c",
   277 => x"04",
   278 => x"42",
   279 => x"98",
   280 => x"60",
   281 => x"f8",
   282 => x"41",
   283 => x"fa",
   284 => x"00",
   285 => x"4e",
   286 => x"21",
   287 => x"c8",
   288 => x"00",
   289 => x"64",
   290 => x"41",
   291 => x"fa",
   292 => x"00",
   293 => x"54",
   294 => x"21",
   295 => x"c8",
   296 => x"00",
   297 => x"68",
   298 => x"41",
   299 => x"fa",
   300 => x"00",
   301 => x"5a",
   302 => x"21",
   303 => x"c8",
   304 => x"00",
   305 => x"6c",
   306 => x"41",
   307 => x"fa",
   308 => x"00",
   309 => x"60",
   310 => x"21",
   311 => x"c8",
   312 => x"00",
   313 => x"70",
   314 => x"41",
   315 => x"fa",
   316 => x"00",
   317 => x"66",
   318 => x"21",
   319 => x"c8",
   320 => x"00",
   321 => x"74",
   322 => x"41",
   323 => x"fa",
   324 => x"00",
   325 => x"6c",
   326 => x"21",
   327 => x"c8",
   328 => x"00",
   329 => x"78",
   330 => x"41",
   331 => x"fa",
   332 => x"00",
   333 => x"72",
   334 => x"21",
   335 => x"c8",
   336 => x"00",
   337 => x"7c",
   338 => x"48",
   339 => x"78",
   340 => x"00",
   341 => x"01",
   342 => x"48",
   343 => x"7a",
   344 => x"00",
   345 => x"0a",
   346 => x"4e",
   347 => x"b9",
   348 => x"00",
   349 => x"00",
   350 => x"02",
   351 => x"80",
   352 => x"60",
   353 => x"fe",
   354 => x"42",
   355 => x"6f",
   356 => x"6f",
   357 => x"74",
   358 => x"72",
   359 => x"6f",
   360 => x"6d",
   361 => x"00",
   362 => x"48",
   363 => x"e7",
   364 => x"ff",
   365 => x"fe",
   366 => x"48",
   367 => x"7a",
   368 => x"00",
   369 => x"5c",
   370 => x"2f",
   371 => x"3a",
   372 => x"00",
   373 => x"60",
   374 => x"4e",
   375 => x"75",
   376 => x"48",
   377 => x"e7",
   378 => x"ff",
   379 => x"fe",
   380 => x"48",
   381 => x"7a",
   382 => x"00",
   383 => x"4e",
   384 => x"2f",
   385 => x"3a",
   386 => x"00",
   387 => x"56",
   388 => x"4e",
   389 => x"75",
   390 => x"48",
   391 => x"e7",
   392 => x"ff",
   393 => x"fe",
   394 => x"48",
   395 => x"7a",
   396 => x"00",
   397 => x"40",
   398 => x"2f",
   399 => x"3a",
   400 => x"00",
   401 => x"4c",
   402 => x"4e",
   403 => x"75",
   404 => x"48",
   405 => x"e7",
   406 => x"ff",
   407 => x"fe",
   408 => x"48",
   409 => x"7a",
   410 => x"00",
   411 => x"32",
   412 => x"2f",
   413 => x"3a",
   414 => x"00",
   415 => x"42",
   416 => x"4e",
   417 => x"75",
   418 => x"48",
   419 => x"e7",
   420 => x"ff",
   421 => x"fe",
   422 => x"48",
   423 => x"7a",
   424 => x"00",
   425 => x"24",
   426 => x"2f",
   427 => x"3a",
   428 => x"00",
   429 => x"38",
   430 => x"4e",
   431 => x"75",
   432 => x"48",
   433 => x"e7",
   434 => x"ff",
   435 => x"fe",
   436 => x"48",
   437 => x"7a",
   438 => x"00",
   439 => x"16",
   440 => x"2f",
   441 => x"3a",
   442 => x"00",
   443 => x"2e",
   444 => x"4e",
   445 => x"75",
   446 => x"48",
   447 => x"e7",
   448 => x"ff",
   449 => x"fe",
   450 => x"48",
   451 => x"7a",
   452 => x"00",
   453 => x"08",
   454 => x"2f",
   455 => x"3a",
   456 => x"00",
   457 => x"24",
   458 => x"4e",
   459 => x"75",
   460 => x"4c",
   461 => x"df",
   462 => x"7f",
   463 => x"ff",
   464 => x"4e",
   465 => x"73",
   466 => x"4e",
   467 => x"75",
   468 => x"00",
   469 => x"00",
   470 => x"01",
   471 => x"d2",
   472 => x"00",
   473 => x"00",
   474 => x"01",
   475 => x"d2",
   476 => x"00",
   477 => x"00",
   478 => x"01",
   479 => x"d2",
   480 => x"00",
   481 => x"00",
   482 => x"01",
   483 => x"d2",
   484 => x"00",
   485 => x"00",
   486 => x"01",
   487 => x"d2",
   488 => x"00",
   489 => x"00",
   490 => x"01",
   491 => x"d2",
   492 => x"00",
   493 => x"00",
   494 => x"01",
   495 => x"d2",
   496 => x"46",
   497 => x"fc",
   498 => x"20",
   499 => x"00",
   500 => x"4e",
   501 => x"75",
   502 => x"46",
   503 => x"fc",
   504 => x"27",
   505 => x"00",
   506 => x"4e",
   507 => x"75",
   508 => x"00",
   509 => x"00",
   510 => x"00",
   511 => x"00",
   512 => x"cf",
   513 => x"00",
   514 => x"00",
   515 => x"00",
   516 => x"00",
   517 => x"00",
   518 => x"00",
   519 => x"00",
   520 => x"8c",
   521 => x"ff",
   522 => x"f0",
   523 => x"00",
   524 => x"00",
   525 => x"00",
   526 => x"00",
   527 => x"00",
   528 => x"08",
   529 => x"cc",
   530 => x"ff",
   531 => x"f0",
   532 => x"00",
   533 => x"00",
   534 => x"00",
   535 => x"00",
   536 => x"08",
   537 => x"cc",
   538 => x"cc",
   539 => x"ff",
   540 => x"ff",
   541 => x"00",
   542 => x"00",
   543 => x"00",
   544 => x"08",
   545 => x"8c",
   546 => x"cc",
   547 => x"cc",
   548 => x"cf",
   549 => x"ff",
   550 => x"00",
   551 => x"00",
   552 => x"00",
   553 => x"8c",
   554 => x"cc",
   555 => x"cc",
   556 => x"cc",
   557 => x"c8",
   558 => x"00",
   559 => x"00",
   560 => x"00",
   561 => x"88",
   562 => x"cc",
   563 => x"cc",
   564 => x"cc",
   565 => x"80",
   566 => x"00",
   567 => x"00",
   568 => x"00",
   569 => x"08",
   570 => x"cc",
   571 => x"cc",
   572 => x"cf",
   573 => x"00",
   574 => x"00",
   575 => x"00",
   576 => x"00",
   577 => x"08",
   578 => x"cc",
   579 => x"cc",
   580 => x"cc",
   581 => x"f0",
   582 => x"00",
   583 => x"00",
   584 => x"00",
   585 => x"08",
   586 => x"8c",
   587 => x"c8",
   588 => x"cc",
   589 => x"cf",
   590 => x"00",
   591 => x"00",
   592 => x"00",
   593 => x"00",
   594 => x"8c",
   595 => x"80",
   596 => x"8c",
   597 => x"cc",
   598 => x"f0",
   599 => x"00",
   600 => x"00",
   601 => x"00",
   602 => x"88",
   603 => x"00",
   604 => x"08",
   605 => x"cc",
   606 => x"cf",
   607 => x"00",
   608 => x"00",
   609 => x"00",
   610 => x"00",
   611 => x"00",
   612 => x"00",
   613 => x"8c",
   614 => x"cc",
   615 => x"f0",
   616 => x"00",
   617 => x"00",
   618 => x"00",
   619 => x"00",
   620 => x"00",
   621 => x"08",
   622 => x"cc",
   623 => x"c8",
   624 => x"00",
   625 => x"00",
   626 => x"00",
   627 => x"00",
   628 => x"00",
   629 => x"00",
   630 => x"8c",
   631 => x"80",
   632 => x"00",
   633 => x"00",
   634 => x"00",
   635 => x"00",
   636 => x"00",
   637 => x"00",
   638 => x"08",
   639 => x"00",
   640 => x"4e",
   641 => x"56",
   642 => x"00",
   643 => x"00",
   644 => x"2f",
   645 => x"0a",
   646 => x"2f",
   647 => x"02",
   648 => x"32",
   649 => x"39",
   650 => x"81",
   651 => x"00",
   652 => x"00",
   653 => x"2a",
   654 => x"02",
   655 => x"81",
   656 => x"00",
   657 => x"00",
   658 => x"ff",
   659 => x"ff",
   660 => x"24",
   661 => x"01",
   662 => x"e5",
   663 => x"8a",
   664 => x"20",
   665 => x"01",
   666 => x"ef",
   667 => x"88",
   668 => x"90",
   669 => x"82",
   670 => x"d2",
   671 => x"80",
   672 => x"e7",
   673 => x"89",
   674 => x"24",
   675 => x"01",
   676 => x"4c",
   677 => x"3c",
   678 => x"2c",
   679 => x"00",
   680 => x"38",
   681 => x"e3",
   682 => x"8e",
   683 => x"39",
   684 => x"e0",
   685 => x"80",
   686 => x"d2",
   687 => x"81",
   688 => x"93",
   689 => x"81",
   690 => x"90",
   691 => x"81",
   692 => x"33",
   693 => x"c0",
   694 => x"81",
   695 => x"00",
   696 => x"00",
   697 => x"02",
   698 => x"48",
   699 => x"79",
   700 => x"00",
   701 => x"00",
   702 => x"0b",
   703 => x"24",
   704 => x"45",
   705 => x"f9",
   706 => x"00",
   707 => x"00",
   708 => x"08",
   709 => x"8a",
   710 => x"4e",
   711 => x"92",
   712 => x"2f",
   713 => x"3c",
   714 => x"00",
   715 => x"01",
   716 => x"00",
   717 => x"00",
   718 => x"4e",
   719 => x"b9",
   720 => x"00",
   721 => x"00",
   722 => x"06",
   723 => x"fe",
   724 => x"50",
   725 => x"8f",
   726 => x"4a",
   727 => x"80",
   728 => x"67",
   729 => x"08",
   730 => x"48",
   731 => x"79",
   732 => x"00",
   733 => x"00",
   734 => x"0b",
   735 => x"41",
   736 => x"60",
   737 => x"06",
   738 => x"48",
   739 => x"79",
   740 => x"00",
   741 => x"00",
   742 => x"0b",
   743 => x"56",
   744 => x"4e",
   745 => x"92",
   746 => x"58",
   747 => x"8f",
   748 => x"42",
   749 => x"80",
   750 => x"24",
   751 => x"2e",
   752 => x"ff",
   753 => x"f8",
   754 => x"24",
   755 => x"6e",
   756 => x"ff",
   757 => x"fc",
   758 => x"4e",
   759 => x"5e",
   760 => x"4e",
   761 => x"75",
   762 => x"00",
   763 => x"00",
   764 => x"4e",
   765 => x"56",
   766 => x"00",
   767 => x"00",
   768 => x"48",
   769 => x"e7",
   770 => x"38",
   771 => x"20",
   772 => x"24",
   773 => x"2e",
   774 => x"00",
   775 => x"08",
   776 => x"67",
   777 => x"3a",
   778 => x"76",
   779 => x"08",
   780 => x"42",
   781 => x"80",
   782 => x"45",
   783 => x"f9",
   784 => x"00",
   785 => x"00",
   786 => x"08",
   787 => x"6c",
   788 => x"22",
   789 => x"02",
   790 => x"78",
   791 => x"1c",
   792 => x"e8",
   793 => x"a9",
   794 => x"20",
   795 => x"41",
   796 => x"e9",
   797 => x"8a",
   798 => x"4a",
   799 => x"81",
   800 => x"67",
   801 => x"0c",
   802 => x"70",
   803 => x"09",
   804 => x"b0",
   805 => x"81",
   806 => x"6c",
   807 => x"0a",
   808 => x"41",
   809 => x"e8",
   810 => x"00",
   811 => x"37",
   812 => x"60",
   813 => x"08",
   814 => x"4a",
   815 => x"80",
   816 => x"67",
   817 => x"0c",
   818 => x"41",
   819 => x"e8",
   820 => x"00",
   821 => x"30",
   822 => x"2f",
   823 => x"08",
   824 => x"4e",
   825 => x"92",
   826 => x"58",
   827 => x"8f",
   828 => x"70",
   829 => x"01",
   830 => x"53",
   831 => x"83",
   832 => x"66",
   833 => x"d2",
   834 => x"60",
   835 => x"0c",
   836 => x"48",
   837 => x"78",
   838 => x"00",
   839 => x"30",
   840 => x"4e",
   841 => x"b9",
   842 => x"00",
   843 => x"00",
   844 => x"08",
   845 => x"6c",
   846 => x"58",
   847 => x"8f",
   848 => x"48",
   849 => x"78",
   850 => x"00",
   851 => x"0a",
   852 => x"4e",
   853 => x"b9",
   854 => x"00",
   855 => x"00",
   856 => x"08",
   857 => x"6c",
   858 => x"42",
   859 => x"80",
   860 => x"4c",
   861 => x"ee",
   862 => x"04",
   863 => x"1c",
   864 => x"ff",
   865 => x"f0",
   866 => x"4e",
   867 => x"5e",
   868 => x"4e",
   869 => x"75",
   870 => x"4e",
   871 => x"56",
   872 => x"00",
   873 => x"00",
   874 => x"20",
   875 => x"6e",
   876 => x"00",
   877 => x"08",
   878 => x"20",
   879 => x"28",
   880 => x"40",
   881 => x"00",
   882 => x"20",
   883 => x"30",
   884 => x"01",
   885 => x"70",
   886 => x"00",
   887 => x"01",
   888 => x"00",
   889 => x"04",
   890 => x"20",
   891 => x"30",
   892 => x"01",
   893 => x"70",
   894 => x"00",
   895 => x"00",
   896 => x"80",
   897 => x"00",
   898 => x"20",
   899 => x"30",
   900 => x"01",
   901 => x"70",
   902 => x"00",
   903 => x"00",
   904 => x"c0",
   905 => x"0c",
   906 => x"20",
   907 => x"30",
   908 => x"01",
   909 => x"70",
   910 => x"00",
   911 => x"00",
   912 => x"c0",
   913 => x"04",
   914 => x"20",
   915 => x"30",
   916 => x"01",
   917 => x"70",
   918 => x"00",
   919 => x"00",
   920 => x"80",
   921 => x"0c",
   922 => x"20",
   923 => x"30",
   924 => x"01",
   925 => x"70",
   926 => x"00",
   927 => x"01",
   928 => x"00",
   929 => x"00",
   930 => x"20",
   931 => x"28",
   932 => x"40",
   933 => x"08",
   934 => x"4e",
   935 => x"5e",
   936 => x"4e",
   937 => x"75",
   938 => x"4e",
   939 => x"56",
   940 => x"00",
   941 => x"00",
   942 => x"48",
   943 => x"e7",
   944 => x"38",
   945 => x"20",
   946 => x"24",
   947 => x"6e",
   948 => x"00",
   949 => x"08",
   950 => x"22",
   951 => x"2e",
   952 => x"00",
   953 => x"0c",
   954 => x"20",
   955 => x"2e",
   956 => x"00",
   957 => x"10",
   958 => x"26",
   959 => x"01",
   960 => x"48",
   961 => x"43",
   962 => x"42",
   963 => x"43",
   964 => x"24",
   965 => x"00",
   966 => x"42",
   967 => x"42",
   968 => x"48",
   969 => x"42",
   970 => x"84",
   971 => x"83",
   972 => x"24",
   973 => x"81",
   974 => x"25",
   975 => x"40",
   976 => x"00",
   977 => x"04",
   978 => x"26",
   979 => x"2a",
   980 => x"00",
   981 => x"02",
   982 => x"b4",
   983 => x"83",
   984 => x"67",
   985 => x"18",
   986 => x"48",
   987 => x"79",
   988 => x"00",
   989 => x"00",
   990 => x"08",
   991 => x"b6",
   992 => x"4e",
   993 => x"b9",
   994 => x"00",
   995 => x"00",
   996 => x"08",
   997 => x"8a",
   998 => x"2f",
   999 => x"03",
  1000 => x"4e",
  1001 => x"ba",
  1002 => x"ff",
  1003 => x"12",
  1004 => x"b5",
  1005 => x"83",
  1006 => x"50",
  1007 => x"8f",
  1008 => x"60",
  1009 => x"02",
  1010 => x"42",
  1011 => x"83",
  1012 => x"48",
  1013 => x"6a",
  1014 => x"00",
  1015 => x"08",
  1016 => x"4e",
  1017 => x"ba",
  1018 => x"ff",
  1019 => x"6c",
  1020 => x"28",
  1021 => x"2a",
  1022 => x"00",
  1023 => x"02",
  1024 => x"58",
  1025 => x"8f",
  1026 => x"b4",
  1027 => x"84",
  1028 => x"67",
  1029 => x"18",
  1030 => x"48",
  1031 => x"79",
  1032 => x"00",
  1033 => x"00",
  1034 => x"08",
  1035 => x"dd",
  1036 => x"4e",
  1037 => x"b9",
  1038 => x"00",
  1039 => x"00",
  1040 => x"08",
  1041 => x"8a",
  1042 => x"2f",
  1043 => x"04",
  1044 => x"4e",
  1045 => x"ba",
  1046 => x"fe",
  1047 => x"e6",
  1048 => x"b9",
  1049 => x"82",
  1050 => x"86",
  1051 => x"82",
  1052 => x"50",
  1053 => x"8f",
  1054 => x"20",
  1055 => x"03",
  1056 => x"4c",
  1057 => x"ee",
  1058 => x"04",
  1059 => x"1c",
  1060 => x"ff",
  1061 => x"f0",
  1062 => x"4e",
  1063 => x"5e",
  1064 => x"4e",
  1065 => x"75",
  1066 => x"4e",
  1067 => x"56",
  1068 => x"00",
  1069 => x"00",
  1070 => x"48",
  1071 => x"e7",
  1072 => x"3f",
  1073 => x"20",
  1074 => x"24",
  1075 => x"6e",
  1076 => x"00",
  1077 => x"08",
  1078 => x"2a",
  1079 => x"2e",
  1080 => x"00",
  1081 => x"0c",
  1082 => x"20",
  1083 => x"2e",
  1084 => x"00",
  1085 => x"10",
  1086 => x"3e",
  1087 => x"00",
  1088 => x"42",
  1089 => x"83",
  1090 => x"36",
  1091 => x"00",
  1092 => x"28",
  1093 => x"05",
  1094 => x"42",
  1095 => x"44",
  1096 => x"88",
  1097 => x"83",
  1098 => x"48",
  1099 => x"43",
  1100 => x"42",
  1101 => x"43",
  1102 => x"86",
  1103 => x"45",
  1104 => x"24",
  1105 => x"85",
  1106 => x"34",
  1107 => x"80",
  1108 => x"24",
  1109 => x"12",
  1110 => x"b6",
  1111 => x"82",
  1112 => x"67",
  1113 => x"18",
  1114 => x"48",
  1115 => x"79",
  1116 => x"00",
  1117 => x"00",
  1118 => x"09",
  1119 => x"04",
  1120 => x"4e",
  1121 => x"b9",
  1122 => x"00",
  1123 => x"00",
  1124 => x"08",
  1125 => x"8a",
  1126 => x"2f",
  1127 => x"02",
  1128 => x"4e",
  1129 => x"ba",
  1130 => x"fe",
  1131 => x"92",
  1132 => x"b7",
  1133 => x"82",
  1134 => x"50",
  1135 => x"8f",
  1136 => x"60",
  1137 => x"02",
  1138 => x"42",
  1139 => x"82",
  1140 => x"2f",
  1141 => x"0a",
  1142 => x"4e",
  1143 => x"ba",
  1144 => x"fe",
  1145 => x"ee",
  1146 => x"2c",
  1147 => x"12",
  1148 => x"58",
  1149 => x"8f",
  1150 => x"b6",
  1151 => x"86",
  1152 => x"67",
  1153 => x"18",
  1154 => x"48",
  1155 => x"79",
  1156 => x"00",
  1157 => x"00",
  1158 => x"09",
  1159 => x"28",
  1160 => x"4e",
  1161 => x"b9",
  1162 => x"00",
  1163 => x"00",
  1164 => x"08",
  1165 => x"8a",
  1166 => x"2f",
  1167 => x"06",
  1168 => x"4e",
  1169 => x"ba",
  1170 => x"fe",
  1171 => x"6a",
  1172 => x"bd",
  1173 => x"83",
  1174 => x"84",
  1175 => x"83",
  1176 => x"50",
  1177 => x"8f",
  1178 => x"25",
  1179 => x"45",
  1180 => x"00",
  1181 => x"04",
  1182 => x"35",
  1183 => x"47",
  1184 => x"00",
  1185 => x"06",
  1186 => x"26",
  1187 => x"2a",
  1188 => x"00",
  1189 => x"04",
  1190 => x"b8",
  1191 => x"83",
  1192 => x"67",
  1193 => x"18",
  1194 => x"48",
  1195 => x"79",
  1196 => x"00",
  1197 => x"00",
  1198 => x"09",
  1199 => x"4c",
  1200 => x"4e",
  1201 => x"b9",
  1202 => x"00",
  1203 => x"00",
  1204 => x"08",
  1205 => x"8a",
  1206 => x"2f",
  1207 => x"03",
  1208 => x"4e",
  1209 => x"ba",
  1210 => x"fe",
  1211 => x"42",
  1212 => x"b9",
  1213 => x"83",
  1214 => x"84",
  1215 => x"83",
  1216 => x"50",
  1217 => x"8f",
  1218 => x"48",
  1219 => x"6a",
  1220 => x"00",
  1221 => x"04",
  1222 => x"4e",
  1223 => x"ba",
  1224 => x"fe",
  1225 => x"9e",
  1226 => x"26",
  1227 => x"2a",
  1228 => x"00",
  1229 => x"04",
  1230 => x"58",
  1231 => x"8f",
  1232 => x"b8",
  1233 => x"83",
  1234 => x"67",
  1235 => x"18",
  1236 => x"48",
  1237 => x"79",
  1238 => x"00",
  1239 => x"00",
  1240 => x"09",
  1241 => x"70",
  1242 => x"4e",
  1243 => x"b9",
  1244 => x"00",
  1245 => x"00",
  1246 => x"08",
  1247 => x"8a",
  1248 => x"2f",
  1249 => x"03",
  1250 => x"4e",
  1251 => x"ba",
  1252 => x"fe",
  1253 => x"18",
  1254 => x"b7",
  1255 => x"84",
  1256 => x"84",
  1257 => x"84",
  1258 => x"50",
  1259 => x"8f",
  1260 => x"20",
  1261 => x"02",
  1262 => x"4c",
  1263 => x"ee",
  1264 => x"04",
  1265 => x"fc",
  1266 => x"ff",
  1267 => x"e4",
  1268 => x"4e",
  1269 => x"5e",
  1270 => x"4e",
  1271 => x"75",
  1272 => x"4e",
  1273 => x"56",
  1274 => x"00",
  1275 => x"00",
  1276 => x"48",
  1277 => x"e7",
  1278 => x"3f",
  1279 => x"3c",
  1280 => x"24",
  1281 => x"6e",
  1282 => x"00",
  1283 => x"08",
  1284 => x"26",
  1285 => x"2e",
  1286 => x"00",
  1287 => x"0c",
  1288 => x"20",
  1289 => x"2e",
  1290 => x"00",
  1291 => x"10",
  1292 => x"42",
  1293 => x"84",
  1294 => x"18",
  1295 => x"00",
  1296 => x"72",
  1297 => x"ff",
  1298 => x"46",
  1299 => x"01",
  1300 => x"c2",
  1301 => x"83",
  1302 => x"82",
  1303 => x"84",
  1304 => x"28",
  1305 => x"41",
  1306 => x"2e",
  1307 => x"04",
  1308 => x"e1",
  1309 => x"8f",
  1310 => x"22",
  1311 => x"03",
  1312 => x"02",
  1313 => x"41",
  1314 => x"00",
  1315 => x"ff",
  1316 => x"8e",
  1317 => x"81",
  1318 => x"2c",
  1319 => x"04",
  1320 => x"48",
  1321 => x"46",
  1322 => x"42",
  1323 => x"46",
  1324 => x"22",
  1325 => x"03",
  1326 => x"02",
  1327 => x"81",
  1328 => x"ff",
  1329 => x"00",
  1330 => x"ff",
  1331 => x"ff",
  1332 => x"8c",
  1333 => x"81",
  1334 => x"2a",
  1335 => x"04",
  1336 => x"72",
  1337 => x"18",
  1338 => x"e3",
  1339 => x"ad",
  1340 => x"22",
  1341 => x"03",
  1342 => x"02",
  1343 => x"81",
  1344 => x"00",
  1345 => x"ff",
  1346 => x"ff",
  1347 => x"ff",
  1348 => x"8a",
  1349 => x"81",
  1350 => x"24",
  1351 => x"83",
  1352 => x"15",
  1353 => x"40",
  1354 => x"00",
  1355 => x"03",
  1356 => x"25",
  1357 => x"43",
  1358 => x"00",
  1359 => x"04",
  1360 => x"15",
  1361 => x"40",
  1362 => x"00",
  1363 => x"06",
  1364 => x"25",
  1365 => x"43",
  1366 => x"00",
  1367 => x"08",
  1368 => x"15",
  1369 => x"40",
  1370 => x"00",
  1371 => x"09",
  1372 => x"25",
  1373 => x"43",
  1374 => x"00",
  1375 => x"0c",
  1376 => x"15",
  1377 => x"40",
  1378 => x"00",
  1379 => x"0c",
  1380 => x"24",
  1381 => x"12",
  1382 => x"b9",
  1383 => x"c2",
  1384 => x"67",
  1385 => x"26",
  1386 => x"48",
  1387 => x"79",
  1388 => x"00",
  1389 => x"00",
  1390 => x"09",
  1391 => x"94",
  1392 => x"4e",
  1393 => x"b9",
  1394 => x"00",
  1395 => x"00",
  1396 => x"08",
  1397 => x"8a",
  1398 => x"2f",
  1399 => x"02",
  1400 => x"47",
  1401 => x"fa",
  1402 => x"fd",
  1403 => x"82",
  1404 => x"4e",
  1405 => x"93",
  1406 => x"2f",
  1407 => x"03",
  1408 => x"4e",
  1409 => x"93",
  1410 => x"2f",
  1411 => x"04",
  1412 => x"4e",
  1413 => x"93",
  1414 => x"20",
  1415 => x"0c",
  1416 => x"b1",
  1417 => x"82",
  1418 => x"4f",
  1419 => x"ef",
  1420 => x"00",
  1421 => x"10",
  1422 => x"60",
  1423 => x"02",
  1424 => x"42",
  1425 => x"82",
  1426 => x"47",
  1427 => x"ea",
  1428 => x"00",
  1429 => x"08",
  1430 => x"2f",
  1431 => x"0b",
  1432 => x"4e",
  1433 => x"ba",
  1434 => x"fd",
  1435 => x"cc",
  1436 => x"2a",
  1437 => x"52",
  1438 => x"58",
  1439 => x"8f",
  1440 => x"b9",
  1441 => x"cd",
  1442 => x"67",
  1443 => x"2a",
  1444 => x"48",
  1445 => x"79",
  1446 => x"00",
  1447 => x"00",
  1448 => x"09",
  1449 => x"b7",
  1450 => x"4e",
  1451 => x"b9",
  1452 => x"00",
  1453 => x"00",
  1454 => x"08",
  1455 => x"8a",
  1456 => x"2f",
  1457 => x"0d",
  1458 => x"4e",
  1459 => x"ba",
  1460 => x"fd",
  1461 => x"48",
  1462 => x"2f",
  1463 => x"03",
  1464 => x"4e",
  1465 => x"ba",
  1466 => x"fd",
  1467 => x"42",
  1468 => x"2f",
  1469 => x"04",
  1470 => x"4e",
  1471 => x"ba",
  1472 => x"fd",
  1473 => x"3c",
  1474 => x"20",
  1475 => x"0c",
  1476 => x"22",
  1477 => x"0d",
  1478 => x"b3",
  1479 => x"80",
  1480 => x"84",
  1481 => x"80",
  1482 => x"4f",
  1483 => x"ef",
  1484 => x"00",
  1485 => x"10",
  1486 => x"28",
  1487 => x"6a",
  1488 => x"00",
  1489 => x"04",
  1490 => x"be",
  1491 => x"8c",
  1492 => x"67",
  1493 => x"26",
  1494 => x"48",
  1495 => x"79",
  1496 => x"00",
  1497 => x"00",
  1498 => x"09",
  1499 => x"da",
  1500 => x"4e",
  1501 => x"b9",
  1502 => x"00",
  1503 => x"00",
  1504 => x"08",
  1505 => x"8a",
  1506 => x"2f",
  1507 => x"0c",
  1508 => x"4b",
  1509 => x"fa",
  1510 => x"fd",
  1511 => x"16",
  1512 => x"4e",
  1513 => x"95",
  1514 => x"2f",
  1515 => x"03",
  1516 => x"4e",
  1517 => x"95",
  1518 => x"2f",
  1519 => x"04",
  1520 => x"4e",
  1521 => x"95",
  1522 => x"20",
  1523 => x"0c",
  1524 => x"bf",
  1525 => x"80",
  1526 => x"84",
  1527 => x"80",
  1528 => x"4f",
  1529 => x"ef",
  1530 => x"00",
  1531 => x"10",
  1532 => x"2f",
  1533 => x"0b",
  1534 => x"4e",
  1535 => x"ba",
  1536 => x"fd",
  1537 => x"66",
  1538 => x"28",
  1539 => x"6a",
  1540 => x"00",
  1541 => x"04",
  1542 => x"58",
  1543 => x"8f",
  1544 => x"be",
  1545 => x"8c",
  1546 => x"67",
  1547 => x"26",
  1548 => x"48",
  1549 => x"79",
  1550 => x"00",
  1551 => x"00",
  1552 => x"09",
  1553 => x"fd",
  1554 => x"4e",
  1555 => x"b9",
  1556 => x"00",
  1557 => x"00",
  1558 => x"08",
  1559 => x"8a",
  1560 => x"2f",
  1561 => x"0c",
  1562 => x"4b",
  1563 => x"fa",
  1564 => x"fc",
  1565 => x"e0",
  1566 => x"4e",
  1567 => x"95",
  1568 => x"2f",
  1569 => x"03",
  1570 => x"4e",
  1571 => x"95",
  1572 => x"2f",
  1573 => x"04",
  1574 => x"4e",
  1575 => x"95",
  1576 => x"20",
  1577 => x"0c",
  1578 => x"b1",
  1579 => x"87",
  1580 => x"84",
  1581 => x"87",
  1582 => x"4f",
  1583 => x"ef",
  1584 => x"00",
  1585 => x"10",
  1586 => x"2e",
  1587 => x"2a",
  1588 => x"00",
  1589 => x"08",
  1590 => x"bc",
  1591 => x"87",
  1592 => x"67",
  1593 => x"24",
  1594 => x"48",
  1595 => x"79",
  1596 => x"00",
  1597 => x"00",
  1598 => x"0a",
  1599 => x"20",
  1600 => x"4e",
  1601 => x"b9",
  1602 => x"00",
  1603 => x"00",
  1604 => x"08",
  1605 => x"8a",
  1606 => x"2f",
  1607 => x"07",
  1608 => x"49",
  1609 => x"fa",
  1610 => x"fc",
  1611 => x"b2",
  1612 => x"4e",
  1613 => x"94",
  1614 => x"2f",
  1615 => x"03",
  1616 => x"4e",
  1617 => x"94",
  1618 => x"2f",
  1619 => x"04",
  1620 => x"4e",
  1621 => x"94",
  1622 => x"bd",
  1623 => x"87",
  1624 => x"84",
  1625 => x"87",
  1626 => x"4f",
  1627 => x"ef",
  1628 => x"00",
  1629 => x"10",
  1630 => x"2f",
  1631 => x"0b",
  1632 => x"4e",
  1633 => x"ba",
  1634 => x"fd",
  1635 => x"04",
  1636 => x"2e",
  1637 => x"2a",
  1638 => x"00",
  1639 => x"08",
  1640 => x"58",
  1641 => x"8f",
  1642 => x"bc",
  1643 => x"87",
  1644 => x"67",
  1645 => x"24",
  1646 => x"48",
  1647 => x"79",
  1648 => x"00",
  1649 => x"00",
  1650 => x"0a",
  1651 => x"43",
  1652 => x"4e",
  1653 => x"b9",
  1654 => x"00",
  1655 => x"00",
  1656 => x"08",
  1657 => x"8a",
  1658 => x"2f",
  1659 => x"07",
  1660 => x"49",
  1661 => x"fa",
  1662 => x"fc",
  1663 => x"7e",
  1664 => x"4e",
  1665 => x"94",
  1666 => x"2f",
  1667 => x"03",
  1668 => x"4e",
  1669 => x"94",
  1670 => x"2f",
  1671 => x"04",
  1672 => x"4e",
  1673 => x"94",
  1674 => x"bf",
  1675 => x"86",
  1676 => x"84",
  1677 => x"86",
  1678 => x"4f",
  1679 => x"ef",
  1680 => x"00",
  1681 => x"10",
  1682 => x"2c",
  1683 => x"2a",
  1684 => x"00",
  1685 => x"0c",
  1686 => x"ba",
  1687 => x"86",
  1688 => x"67",
  1689 => x"24",
  1690 => x"48",
  1691 => x"79",
  1692 => x"00",
  1693 => x"00",
  1694 => x"0a",
  1695 => x"66",
  1696 => x"4e",
  1697 => x"b9",
  1698 => x"00",
  1699 => x"00",
  1700 => x"08",
  1701 => x"8a",
  1702 => x"2f",
  1703 => x"06",
  1704 => x"49",
  1705 => x"fa",
  1706 => x"fc",
  1707 => x"52",
  1708 => x"4e",
  1709 => x"94",
  1710 => x"2f",
  1711 => x"03",
  1712 => x"4e",
  1713 => x"94",
  1714 => x"2f",
  1715 => x"04",
  1716 => x"4e",
  1717 => x"94",
  1718 => x"bb",
  1719 => x"86",
  1720 => x"84",
  1721 => x"86",
  1722 => x"4f",
  1723 => x"ef",
  1724 => x"00",
  1725 => x"10",
  1726 => x"2f",
  1727 => x"0b",
  1728 => x"4e",
  1729 => x"ba",
  1730 => x"fc",
  1731 => x"a4",
  1732 => x"2c",
  1733 => x"2a",
  1734 => x"00",
  1735 => x"0c",
  1736 => x"58",
  1737 => x"8f",
  1738 => x"ba",
  1739 => x"86",
  1740 => x"67",
  1741 => x"24",
  1742 => x"48",
  1743 => x"79",
  1744 => x"00",
  1745 => x"00",
  1746 => x"0a",
  1747 => x"89",
  1748 => x"4e",
  1749 => x"b9",
  1750 => x"00",
  1751 => x"00",
  1752 => x"08",
  1753 => x"8a",
  1754 => x"2f",
  1755 => x"06",
  1756 => x"45",
  1757 => x"fa",
  1758 => x"fc",
  1759 => x"1e",
  1760 => x"4e",
  1761 => x"92",
  1762 => x"2f",
  1763 => x"03",
  1764 => x"4e",
  1765 => x"92",
  1766 => x"2f",
  1767 => x"04",
  1768 => x"4e",
  1769 => x"92",
  1770 => x"bd",
  1771 => x"85",
  1772 => x"84",
  1773 => x"85",
  1774 => x"4f",
  1775 => x"ef",
  1776 => x"00",
  1777 => x"10",
  1778 => x"20",
  1779 => x"02",
  1780 => x"4c",
  1781 => x"ee",
  1782 => x"3c",
  1783 => x"fc",
  1784 => x"ff",
  1785 => x"d8",
  1786 => x"4e",
  1787 => x"5e",
  1788 => x"4e",
  1789 => x"75",
  1790 => x"4e",
  1791 => x"56",
  1792 => x"00",
  1793 => x"00",
  1794 => x"48",
  1795 => x"e7",
  1796 => x"3f",
  1797 => x"30",
  1798 => x"2e",
  1799 => x"2e",
  1800 => x"00",
  1801 => x"08",
  1802 => x"48",
  1803 => x"79",
  1804 => x"00",
  1805 => x"00",
  1806 => x"0a",
  1807 => x"ac",
  1808 => x"4e",
  1809 => x"b9",
  1810 => x"00",
  1811 => x"00",
  1812 => x"08",
  1813 => x"8a",
  1814 => x"58",
  1815 => x"8f",
  1816 => x"42",
  1817 => x"83",
  1818 => x"42",
  1819 => x"82",
  1820 => x"47",
  1821 => x"fa",
  1822 => x"fd",
  1823 => x"0c",
  1824 => x"45",
  1825 => x"f9",
  1826 => x"00",
  1827 => x"00",
  1828 => x"08",
  1829 => x"6c",
  1830 => x"60",
  1831 => x"34",
  1832 => x"3f",
  1833 => x"04",
  1834 => x"42",
  1835 => x"67",
  1836 => x"2f",
  1837 => x"03",
  1838 => x"2f",
  1839 => x"07",
  1840 => x"4e",
  1841 => x"93",
  1842 => x"84",
  1843 => x"80",
  1844 => x"06",
  1845 => x"84",
  1846 => x"00",
  1847 => x"31",
  1848 => x"87",
  1849 => x"65",
  1850 => x"4f",
  1851 => x"ef",
  1852 => x"00",
  1853 => x"0c",
  1854 => x"0c",
  1855 => x"84",
  1856 => x"80",
  1857 => x"14",
  1858 => x"1f",
  1859 => x"2e",
  1860 => x"66",
  1861 => x"e2",
  1862 => x"48",
  1863 => x"78",
  1864 => x"00",
  1865 => x"2e",
  1866 => x"4e",
  1867 => x"92",
  1868 => x"06",
  1869 => x"83",
  1870 => x"00",
  1871 => x"21",
  1872 => x"23",
  1873 => x"45",
  1874 => x"58",
  1875 => x"8f",
  1876 => x"0c",
  1877 => x"83",
  1878 => x"80",
  1879 => x"05",
  1880 => x"41",
  1881 => x"91",
  1882 => x"67",
  1883 => x"04",
  1884 => x"42",
  1885 => x"84",
  1886 => x"60",
  1887 => x"c8",
  1888 => x"4a",
  1889 => x"82",
  1890 => x"67",
  1891 => x"18",
  1892 => x"48",
  1893 => x"79",
  1894 => x"00",
  1895 => x"00",
  1896 => x"0a",
  1897 => x"c1",
  1898 => x"4e",
  1899 => x"b9",
  1900 => x"00",
  1901 => x"00",
  1902 => x"08",
  1903 => x"8a",
  1904 => x"2f",
  1905 => x"02",
  1906 => x"4e",
  1907 => x"ba",
  1908 => x"fb",
  1909 => x"88",
  1910 => x"50",
  1911 => x"8f",
  1912 => x"42",
  1913 => x"84",
  1914 => x"60",
  1915 => x"02",
  1916 => x"78",
  1917 => x"01",
  1918 => x"48",
  1919 => x"79",
  1920 => x"00",
  1921 => x"00",
  1922 => x"0a",
  1923 => x"e1",
  1924 => x"4e",
  1925 => x"b9",
  1926 => x"00",
  1927 => x"00",
  1928 => x"08",
  1929 => x"8a",
  1930 => x"58",
  1931 => x"8f",
  1932 => x"42",
  1933 => x"85",
  1934 => x"42",
  1935 => x"83",
  1936 => x"47",
  1937 => x"fa",
  1938 => x"fc",
  1939 => x"18",
  1940 => x"45",
  1941 => x"f9",
  1942 => x"00",
  1943 => x"00",
  1944 => x"08",
  1945 => x"6c",
  1946 => x"60",
  1947 => x"32",
  1948 => x"2f",
  1949 => x"06",
  1950 => x"2f",
  1951 => x"05",
  1952 => x"2f",
  1953 => x"07",
  1954 => x"4e",
  1955 => x"93",
  1956 => x"86",
  1957 => x"80",
  1958 => x"06",
  1959 => x"86",
  1960 => x"00",
  1961 => x"19",
  1962 => x"87",
  1963 => x"65",
  1964 => x"4f",
  1965 => x"ef",
  1966 => x"00",
  1967 => x"0c",
  1968 => x"0c",
  1969 => x"86",
  1970 => x"80",
  1971 => x"0b",
  1972 => x"16",
  1973 => x"94",
  1974 => x"66",
  1975 => x"e4",
  1976 => x"48",
  1977 => x"78",
  1978 => x"00",
  1979 => x"2e",
  1980 => x"4e",
  1981 => x"92",
  1982 => x"06",
  1983 => x"85",
  1984 => x"00",
  1985 => x"13",
  1986 => x"45",
  1987 => x"67",
  1988 => x"58",
  1989 => x"8f",
  1990 => x"0c",
  1991 => x"85",
  1992 => x"80",
  1993 => x"0c",
  1994 => x"25",
  1995 => x"63",
  1996 => x"67",
  1997 => x"04",
  1998 => x"42",
  1999 => x"86",
  2000 => x"60",
  2001 => x"ca",
  2002 => x"4a",
  2003 => x"83",
  2004 => x"67",
  2005 => x"0a",
  2006 => x"2f",
  2007 => x"03",
  2008 => x"4e",
  2009 => x"ba",
  2010 => x"fb",
  2011 => x"22",
  2012 => x"58",
  2013 => x"8f",
  2014 => x"42",
  2015 => x"84",
  2016 => x"86",
  2017 => x"82",
  2018 => x"48",
  2019 => x"79",
  2020 => x"00",
  2021 => x"00",
  2022 => x"0a",
  2023 => x"fb",
  2024 => x"4e",
  2025 => x"b9",
  2026 => x"00",
  2027 => x"00",
  2028 => x"08",
  2029 => x"8a",
  2030 => x"58",
  2031 => x"8f",
  2032 => x"42",
  2033 => x"85",
  2034 => x"42",
  2035 => x"82",
  2036 => x"47",
  2037 => x"fa",
  2038 => x"fd",
  2039 => x"02",
  2040 => x"45",
  2041 => x"f9",
  2042 => x"00",
  2043 => x"00",
  2044 => x"08",
  2045 => x"6c",
  2046 => x"60",
  2047 => x"36",
  2048 => x"42",
  2049 => x"80",
  2050 => x"10",
  2051 => x"06",
  2052 => x"2f",
  2053 => x"00",
  2054 => x"2f",
  2055 => x"05",
  2056 => x"2f",
  2057 => x"07",
  2058 => x"4e",
  2059 => x"93",
  2060 => x"84",
  2061 => x"80",
  2062 => x"06",
  2063 => x"86",
  2064 => x"00",
  2065 => x"28",
  2066 => x"76",
  2067 => x"53",
  2068 => x"4f",
  2069 => x"ef",
  2070 => x"00",
  2071 => x"0c",
  2072 => x"0c",
  2073 => x"86",
  2074 => x"80",
  2075 => x"06",
  2076 => x"62",
  2077 => x"9e",
  2078 => x"66",
  2079 => x"e0",
  2080 => x"48",
  2081 => x"78",
  2082 => x"00",
  2083 => x"2e",
  2084 => x"4e",
  2085 => x"92",
  2086 => x"06",
  2087 => x"85",
  2088 => x"00",
  2089 => x"71",
  2090 => x"23",
  2091 => x"41",
  2092 => x"58",
  2093 => x"8f",
  2094 => x"0c",
  2095 => x"85",
  2096 => x"80",
  2097 => x"29",
  2098 => x"ef",
  2099 => x"a2",
  2100 => x"67",
  2101 => x"04",
  2102 => x"42",
  2103 => x"86",
  2104 => x"60",
  2105 => x"c6",
  2106 => x"4a",
  2107 => x"82",
  2108 => x"67",
  2109 => x"0a",
  2110 => x"2f",
  2111 => x"02",
  2112 => x"4e",
  2113 => x"ba",
  2114 => x"fa",
  2115 => x"ba",
  2116 => x"58",
  2117 => x"8f",
  2118 => x"42",
  2119 => x"84",
  2120 => x"84",
  2121 => x"83",
  2122 => x"67",
  2123 => x"14",
  2124 => x"48",
  2125 => x"79",
  2126 => x"00",
  2127 => x"00",
  2128 => x"0b",
  2129 => x"10",
  2130 => x"4e",
  2131 => x"b9",
  2132 => x"00",
  2133 => x"00",
  2134 => x"08",
  2135 => x"8a",
  2136 => x"2f",
  2137 => x"02",
  2138 => x"4e",
  2139 => x"ba",
  2140 => x"fa",
  2141 => x"a0",
  2142 => x"50",
  2143 => x"8f",
  2144 => x"20",
  2145 => x"04",
  2146 => x"4c",
  2147 => x"ee",
  2148 => x"0c",
  2149 => x"fc",
  2150 => x"ff",
  2151 => x"e0",
  2152 => x"4e",
  2153 => x"5e",
  2154 => x"4e",
  2155 => x"75",
  2156 => x"4e",
  2157 => x"56",
  2158 => x"00",
  2159 => x"00",
  2160 => x"20",
  2161 => x"2e",
  2162 => x"00",
  2163 => x"08",
  2164 => x"32",
  2165 => x"39",
  2166 => x"81",
  2167 => x"00",
  2168 => x"00",
  2169 => x"00",
  2170 => x"08",
  2171 => x"01",
  2172 => x"00",
  2173 => x"08",
  2174 => x"67",
  2175 => x"f4",
  2176 => x"33",
  2177 => x"c0",
  2178 => x"81",
  2179 => x"00",
  2180 => x"00",
  2181 => x"00",
  2182 => x"4e",
  2183 => x"5e",
  2184 => x"4e",
  2185 => x"75",
  2186 => x"4e",
  2187 => x"56",
  2188 => x"00",
  2189 => x"00",
  2190 => x"48",
  2191 => x"e7",
  2192 => x"20",
  2193 => x"30",
  2194 => x"24",
  2195 => x"6e",
  2196 => x"00",
  2197 => x"08",
  2198 => x"47",
  2199 => x"fa",
  2200 => x"ff",
  2201 => x"d4",
  2202 => x"60",
  2203 => x"0a",
  2204 => x"49",
  2205 => x"c0",
  2206 => x"2f",
  2207 => x"00",
  2208 => x"4e",
  2209 => x"93",
  2210 => x"52",
  2211 => x"82",
  2212 => x"58",
  2213 => x"8f",
  2214 => x"10",
  2215 => x"1a",
  2216 => x"66",
  2217 => x"f2",
  2218 => x"20",
  2219 => x"02",
  2220 => x"4c",
  2221 => x"ee",
  2222 => x"0c",
  2223 => x"04",
  2224 => x"ff",
  2225 => x"f4",
  2226 => x"4e",
  2227 => x"5e",
  2228 => x"4e",
  2229 => x"75",
  2230 => x"4d",
  2231 => x"69",
  2232 => x"73",
  2233 => x"61",
  2234 => x"6c",
  2235 => x"69",
  2236 => x"67",
  2237 => x"6e",
  2238 => x"65",
  2239 => x"64",
  2240 => x"20",
  2241 => x"6c",
  2242 => x"6f",
  2243 => x"6e",
  2244 => x"67",
  2245 => x"20",
  2246 => x"63",
  2247 => x"68",
  2248 => x"65",
  2249 => x"63",
  2250 => x"6b",
  2251 => x"20",
  2252 => x"28",
  2253 => x"63",
  2254 => x"61",
  2255 => x"63",
  2256 => x"68",
  2257 => x"65",
  2258 => x"29",
  2259 => x"20",
  2260 => x"66",
  2261 => x"61",
  2262 => x"69",
  2263 => x"6c",
  2264 => x"65",
  2265 => x"64",
  2266 => x"3a",
  2267 => x"20",
  2268 => x"00",
  2269 => x"4d",
  2270 => x"69",
  2271 => x"73",
  2272 => x"61",
  2273 => x"6c",
  2274 => x"69",
  2275 => x"67",
  2276 => x"6e",
  2277 => x"65",
  2278 => x"64",
  2279 => x"20",
  2280 => x"6c",
  2281 => x"6f",
  2282 => x"6e",
  2283 => x"67",
  2284 => x"20",
  2285 => x"63",
  2286 => x"68",
  2287 => x"65",
  2288 => x"63",
  2289 => x"6b",
  2290 => x"20",
  2291 => x"28",
  2292 => x"66",
  2293 => x"6c",
  2294 => x"75",
  2295 => x"73",
  2296 => x"68",
  2297 => x"29",
  2298 => x"20",
  2299 => x"66",
  2300 => x"61",
  2301 => x"69",
  2302 => x"6c",
  2303 => x"65",
  2304 => x"64",
  2305 => x"3a",
  2306 => x"20",
  2307 => x"00",
  2308 => x"4c",
  2309 => x"6f",
  2310 => x"6e",
  2311 => x"67",
  2312 => x"20",
  2313 => x"53",
  2314 => x"68",
  2315 => x"6f",
  2316 => x"72",
  2317 => x"74",
  2318 => x"20",
  2319 => x"63",
  2320 => x"68",
  2321 => x"65",
  2322 => x"63",
  2323 => x"6b",
  2324 => x"20",
  2325 => x"31",
  2326 => x"20",
  2327 => x"28",
  2328 => x"63",
  2329 => x"61",
  2330 => x"63",
  2331 => x"68",
  2332 => x"65",
  2333 => x"29",
  2334 => x"20",
  2335 => x"66",
  2336 => x"61",
  2337 => x"69",
  2338 => x"6c",
  2339 => x"65",
  2340 => x"64",
  2341 => x"3a",
  2342 => x"20",
  2343 => x"00",
  2344 => x"4c",
  2345 => x"6f",
  2346 => x"6e",
  2347 => x"67",
  2348 => x"20",
  2349 => x"53",
  2350 => x"68",
  2351 => x"6f",
  2352 => x"72",
  2353 => x"74",
  2354 => x"20",
  2355 => x"63",
  2356 => x"68",
  2357 => x"65",
  2358 => x"63",
  2359 => x"6b",
  2360 => x"20",
  2361 => x"31",
  2362 => x"20",
  2363 => x"28",
  2364 => x"66",
  2365 => x"6c",
  2366 => x"75",
  2367 => x"73",
  2368 => x"68",
  2369 => x"29",
  2370 => x"20",
  2371 => x"66",
  2372 => x"61",
  2373 => x"69",
  2374 => x"6c",
  2375 => x"65",
  2376 => x"64",
  2377 => x"3a",
  2378 => x"20",
  2379 => x"00",
  2380 => x"4c",
  2381 => x"6f",
  2382 => x"6e",
  2383 => x"67",
  2384 => x"20",
  2385 => x"53",
  2386 => x"68",
  2387 => x"6f",
  2388 => x"72",
  2389 => x"74",
  2390 => x"20",
  2391 => x"63",
  2392 => x"68",
  2393 => x"65",
  2394 => x"63",
  2395 => x"6b",
  2396 => x"20",
  2397 => x"32",
  2398 => x"20",
  2399 => x"28",
  2400 => x"63",
  2401 => x"61",
  2402 => x"63",
  2403 => x"68",
  2404 => x"65",
  2405 => x"29",
  2406 => x"20",
  2407 => x"66",
  2408 => x"61",
  2409 => x"69",
  2410 => x"6c",
  2411 => x"65",
  2412 => x"64",
  2413 => x"3a",
  2414 => x"20",
  2415 => x"00",
  2416 => x"4c",
  2417 => x"6f",
  2418 => x"6e",
  2419 => x"67",
  2420 => x"20",
  2421 => x"53",
  2422 => x"68",
  2423 => x"6f",
  2424 => x"72",
  2425 => x"74",
  2426 => x"20",
  2427 => x"63",
  2428 => x"68",
  2429 => x"65",
  2430 => x"63",
  2431 => x"6b",
  2432 => x"20",
  2433 => x"32",
  2434 => x"20",
  2435 => x"28",
  2436 => x"66",
  2437 => x"6c",
  2438 => x"75",
  2439 => x"73",
  2440 => x"68",
  2441 => x"29",
  2442 => x"20",
  2443 => x"66",
  2444 => x"61",
  2445 => x"69",
  2446 => x"6c",
  2447 => x"65",
  2448 => x"64",
  2449 => x"3a",
  2450 => x"20",
  2451 => x"00",
  2452 => x"4c",
  2453 => x"6f",
  2454 => x"6e",
  2455 => x"67",
  2456 => x"20",
  2457 => x"42",
  2458 => x"79",
  2459 => x"74",
  2460 => x"65",
  2461 => x"20",
  2462 => x"63",
  2463 => x"68",
  2464 => x"65",
  2465 => x"63",
  2466 => x"6b",
  2467 => x"20",
  2468 => x"31",
  2469 => x"20",
  2470 => x"28",
  2471 => x"63",
  2472 => x"61",
  2473 => x"63",
  2474 => x"68",
  2475 => x"65",
  2476 => x"29",
  2477 => x"20",
  2478 => x"66",
  2479 => x"61",
  2480 => x"69",
  2481 => x"6c",
  2482 => x"65",
  2483 => x"64",
  2484 => x"3a",
  2485 => x"20",
  2486 => x"00",
  2487 => x"4c",
  2488 => x"6f",
  2489 => x"6e",
  2490 => x"67",
  2491 => x"20",
  2492 => x"42",
  2493 => x"79",
  2494 => x"74",
  2495 => x"65",
  2496 => x"20",
  2497 => x"63",
  2498 => x"68",
  2499 => x"65",
  2500 => x"63",
  2501 => x"6b",
  2502 => x"20",
  2503 => x"31",
  2504 => x"20",
  2505 => x"28",
  2506 => x"66",
  2507 => x"6c",
  2508 => x"75",
  2509 => x"73",
  2510 => x"68",
  2511 => x"29",
  2512 => x"20",
  2513 => x"66",
  2514 => x"61",
  2515 => x"69",
  2516 => x"6c",
  2517 => x"65",
  2518 => x"64",
  2519 => x"3a",
  2520 => x"20",
  2521 => x"00",
  2522 => x"4c",
  2523 => x"6f",
  2524 => x"6e",
  2525 => x"67",
  2526 => x"20",
  2527 => x"42",
  2528 => x"79",
  2529 => x"74",
  2530 => x"65",
  2531 => x"20",
  2532 => x"63",
  2533 => x"68",
  2534 => x"65",
  2535 => x"63",
  2536 => x"6b",
  2537 => x"20",
  2538 => x"32",
  2539 => x"20",
  2540 => x"28",
  2541 => x"63",
  2542 => x"61",
  2543 => x"63",
  2544 => x"68",
  2545 => x"65",
  2546 => x"29",
  2547 => x"20",
  2548 => x"66",
  2549 => x"61",
  2550 => x"69",
  2551 => x"6c",
  2552 => x"65",
  2553 => x"64",
  2554 => x"3a",
  2555 => x"20",
  2556 => x"00",
  2557 => x"4c",
  2558 => x"6f",
  2559 => x"6e",
  2560 => x"67",
  2561 => x"20",
  2562 => x"42",
  2563 => x"79",
  2564 => x"74",
  2565 => x"65",
  2566 => x"20",
  2567 => x"63",
  2568 => x"68",
  2569 => x"65",
  2570 => x"63",
  2571 => x"6b",
  2572 => x"20",
  2573 => x"32",
  2574 => x"20",
  2575 => x"28",
  2576 => x"66",
  2577 => x"6c",
  2578 => x"75",
  2579 => x"73",
  2580 => x"68",
  2581 => x"29",
  2582 => x"20",
  2583 => x"66",
  2584 => x"61",
  2585 => x"69",
  2586 => x"6c",
  2587 => x"65",
  2588 => x"64",
  2589 => x"3a",
  2590 => x"20",
  2591 => x"00",
  2592 => x"4c",
  2593 => x"6f",
  2594 => x"6e",
  2595 => x"67",
  2596 => x"20",
  2597 => x"42",
  2598 => x"79",
  2599 => x"74",
  2600 => x"65",
  2601 => x"20",
  2602 => x"63",
  2603 => x"68",
  2604 => x"65",
  2605 => x"63",
  2606 => x"6b",
  2607 => x"20",
  2608 => x"33",
  2609 => x"20",
  2610 => x"28",
  2611 => x"63",
  2612 => x"61",
  2613 => x"63",
  2614 => x"68",
  2615 => x"65",
  2616 => x"29",
  2617 => x"20",
  2618 => x"66",
  2619 => x"61",
  2620 => x"69",
  2621 => x"6c",
  2622 => x"65",
  2623 => x"64",
  2624 => x"3a",
  2625 => x"20",
  2626 => x"00",
  2627 => x"4c",
  2628 => x"6f",
  2629 => x"6e",
  2630 => x"67",
  2631 => x"20",
  2632 => x"42",
  2633 => x"79",
  2634 => x"74",
  2635 => x"65",
  2636 => x"20",
  2637 => x"63",
  2638 => x"68",
  2639 => x"65",
  2640 => x"63",
  2641 => x"6b",
  2642 => x"20",
  2643 => x"33",
  2644 => x"20",
  2645 => x"28",
  2646 => x"66",
  2647 => x"6c",
  2648 => x"75",
  2649 => x"73",
  2650 => x"68",
  2651 => x"29",
  2652 => x"20",
  2653 => x"66",
  2654 => x"61",
  2655 => x"69",
  2656 => x"6c",
  2657 => x"65",
  2658 => x"64",
  2659 => x"3a",
  2660 => x"20",
  2661 => x"00",
  2662 => x"4c",
  2663 => x"6f",
  2664 => x"6e",
  2665 => x"67",
  2666 => x"20",
  2667 => x"42",
  2668 => x"79",
  2669 => x"74",
  2670 => x"65",
  2671 => x"20",
  2672 => x"63",
  2673 => x"68",
  2674 => x"65",
  2675 => x"63",
  2676 => x"6b",
  2677 => x"20",
  2678 => x"34",
  2679 => x"20",
  2680 => x"28",
  2681 => x"63",
  2682 => x"61",
  2683 => x"63",
  2684 => x"68",
  2685 => x"65",
  2686 => x"29",
  2687 => x"20",
  2688 => x"66",
  2689 => x"61",
  2690 => x"69",
  2691 => x"6c",
  2692 => x"65",
  2693 => x"64",
  2694 => x"3a",
  2695 => x"20",
  2696 => x"00",
  2697 => x"4c",
  2698 => x"6f",
  2699 => x"6e",
  2700 => x"67",
  2701 => x"20",
  2702 => x"42",
  2703 => x"79",
  2704 => x"74",
  2705 => x"65",
  2706 => x"20",
  2707 => x"63",
  2708 => x"68",
  2709 => x"65",
  2710 => x"63",
  2711 => x"6b",
  2712 => x"20",
  2713 => x"34",
  2714 => x"20",
  2715 => x"28",
  2716 => x"66",
  2717 => x"6c",
  2718 => x"75",
  2719 => x"73",
  2720 => x"68",
  2721 => x"29",
  2722 => x"20",
  2723 => x"66",
  2724 => x"61",
  2725 => x"69",
  2726 => x"6c",
  2727 => x"65",
  2728 => x"64",
  2729 => x"3a",
  2730 => x"20",
  2731 => x"00",
  2732 => x"0a",
  2733 => x"4c",
  2734 => x"6f",
  2735 => x"6e",
  2736 => x"67",
  2737 => x"2f",
  2738 => x"73",
  2739 => x"68",
  2740 => x"6f",
  2741 => x"72",
  2742 => x"74",
  2743 => x"20",
  2744 => x"74",
  2745 => x"65",
  2746 => x"73",
  2747 => x"74",
  2748 => x"2e",
  2749 => x"2e",
  2750 => x"2e",
  2751 => x"0a",
  2752 => x"00",
  2753 => x"42",
  2754 => x"61",
  2755 => x"64",
  2756 => x"20",
  2757 => x"62",
  2758 => x"69",
  2759 => x"74",
  2760 => x"73",
  2761 => x"20",
  2762 => x"66",
  2763 => x"72",
  2764 => x"6f",
  2765 => x"6d",
  2766 => x"20",
  2767 => x"4c",
  2768 => x"6f",
  2769 => x"6e",
  2770 => x"67",
  2771 => x"20",
  2772 => x"53",
  2773 => x"68",
  2774 => x"6f",
  2775 => x"72",
  2776 => x"74",
  2777 => x"20",
  2778 => x"74",
  2779 => x"65",
  2780 => x"73",
  2781 => x"74",
  2782 => x"3a",
  2783 => x"20",
  2784 => x"00",
  2785 => x"0a",
  2786 => x"4d",
  2787 => x"69",
  2788 => x"73",
  2789 => x"61",
  2790 => x"6c",
  2791 => x"69",
  2792 => x"67",
  2793 => x"6e",
  2794 => x"65",
  2795 => x"64",
  2796 => x"20",
  2797 => x"4c",
  2798 => x"6f",
  2799 => x"6e",
  2800 => x"67",
  2801 => x"20",
  2802 => x"74",
  2803 => x"65",
  2804 => x"73",
  2805 => x"74",
  2806 => x"2e",
  2807 => x"2e",
  2808 => x"2e",
  2809 => x"0a",
  2810 => x"00",
  2811 => x"4c",
  2812 => x"6f",
  2813 => x"6e",
  2814 => x"67",
  2815 => x"20",
  2816 => x"2f",
  2817 => x"20",
  2818 => x"62",
  2819 => x"79",
  2820 => x"74",
  2821 => x"65",
  2822 => x"20",
  2823 => x"74",
  2824 => x"65",
  2825 => x"73",
  2826 => x"74",
  2827 => x"2e",
  2828 => x"2e",
  2829 => x"2e",
  2830 => x"0a",
  2831 => x"00",
  2832 => x"42",
  2833 => x"61",
  2834 => x"64",
  2835 => x"20",
  2836 => x"62",
  2837 => x"69",
  2838 => x"74",
  2839 => x"73",
  2840 => x"20",
  2841 => x"64",
  2842 => x"65",
  2843 => x"74",
  2844 => x"65",
  2845 => x"63",
  2846 => x"74",
  2847 => x"65",
  2848 => x"64",
  2849 => x"3a",
  2850 => x"20",
  2851 => x"00",
  2852 => x"43",
  2853 => x"6f",
  2854 => x"6d",
  2855 => x"6d",
  2856 => x"65",
  2857 => x"6e",
  2858 => x"63",
  2859 => x"69",
  2860 => x"6e",
  2861 => x"67",
  2862 => x"20",
  2863 => x"73",
  2864 => x"61",
  2865 => x"6e",
  2866 => x"69",
  2867 => x"74",
  2868 => x"79",
  2869 => x"20",
  2870 => x"63",
  2871 => x"68",
  2872 => x"65",
  2873 => x"63",
  2874 => x"6b",
  2875 => x"73",
  2876 => x"2e",
  2877 => x"2e",
  2878 => x"2e",
  2879 => x"0a",
  2880 => x"00",
  2881 => x"4d",
  2882 => x"65",
  2883 => x"6d",
  2884 => x"6f",
  2885 => x"72",
  2886 => x"79",
  2887 => x"20",
  2888 => x"63",
  2889 => x"68",
  2890 => x"65",
  2891 => x"63",
  2892 => x"6b",
  2893 => x"20",
  2894 => x"70",
  2895 => x"61",
  2896 => x"73",
  2897 => x"73",
  2898 => x"65",
  2899 => x"64",
  2900 => x"0a",
  2901 => x"00",
  2902 => x"4d",
  2903 => x"65",
  2904 => x"6d",
  2905 => x"6f",
  2906 => x"72",
  2907 => x"79",
  2908 => x"20",
  2909 => x"63",
  2910 => x"68",
  2911 => x"65",
  2912 => x"63",
  2913 => x"6b",
  2914 => x"20",
  2915 => x"66",
  2916 => x"61",
  2917 => x"69",
  2918 => x"6c",
  2919 => x"65",
  2920 => x"64",
  2921 => x"0a",
  2922 => x"00",
  2923 => x"00",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;

-- VGA controller
-- a module to handle VGA output

-- Self-contained, must generate timings
-- Programmable, must provide hardware registers that will respond to
-- writes.  Registers will include:  (Decode a 4k chunk)

-- 0 / 2   Framebuffer Address - hi and low
--     4   Even row modulo
--     6   Odd row modulo (allows scandoubling)

--     8  HTotal
--     A  HSize (typically 640)
--     C  HBStart
--     E  HBStop

--    10  VTotal
--    12  VSize (typically 480)
--    14  VBStart
--    16  VBStop

--    18  Control:
--     0  Visible
--     1  Resolution - high, low  - alternatively could make pixel clock programmable...
--     7  Character overlay on/off

--   Character buffer (2048 bytes)


-- Present the following signals to the SOC:
--	clk : in std_logic;
--	reset : in std_logic;

--	reg_addr_in : in std_logic_vector(10 downto 0);
--	reg_rw : std_logic;
--	reg_uds : std_logic;	-- only affects char buffer
--	reg_lds : std_logic;

	--		reqin : in std_logic;  -- now generated by VGA module
	--		data_out : out std_logic_vector(15 downto 0); -- now used internally

--		newframe : in std_logic; -- 
--		addrout : buffer std_logic_vector(23 downto 0); -- to SDRAM
--		data_in : in std_logic_vector(15 downto 0);	-- from SDRAM
--		fill : in std_logic; -- High when data is being written from SDRAM controller
--		req : buffer std_logic -- Request service from SDRAM controller

--		hsync : std_logic -- to monitor
--		vsync : std_logic -- to monitor
--		red : std_logic_vector(4 downto 0);		-- 16-bit 5-6-5 output
--		green : std_logic_vector(5 downto 0);
--		blue : std_logic_vector(4 downto 0);




entity vga_controller is
  port (
		clk : in std_logic;
		reset : in std_logic;

		reg_addr_in : in std_logic_vector(11 downto 0); -- from host CPU
		reg_data_in: in std_logic_vector(15 downto 0);
		reg_data_out: out std_logic_vector(15 downto 0);
		reg_rw : in std_logic;
		reg_uds : in std_logic;
		reg_lds : in std_logic;
		reg_dtack : out std_logic;	-- Needed for char ram access.
		reg_req : in std_logic;

		sdr_addrout : buffer std_logic_vector(23 downto 0); -- to SDRAM
		sdr_datain : in std_logic_vector(15 downto 0);	-- from SDRAM
		sdr_fill : in std_logic; -- High when data is being written from SDRAM controller
		sdr_req : buffer std_logic; -- Request service from SDRAM controller
		sdr_reservebank : buffer std_logic; -- Indicate to SDR controller when requests are not critical timewise
		sdr_reserveaddr : buffer std_logic_vector(23 downto 0); -- Indicate to SDR controller when requests are not critical timewise
		sdr_refresh : out std_logic;

		vblank_int : out std_logic;
		hsync : out std_logic; -- to monitor
		vsync : buffer std_logic; -- to monitor
		red : out unsigned(3 downto 0);		-- 16-bit 5-6-5 output
		green : out unsigned(3 downto 0);
		blue : out unsigned(3 downto 0)
	);
end entity;
	
architecture rtl of vga_controller is
	signal vga_pointer : std_logic_vector(23 downto 0);

	signal framebuffer_pointer : std_logic_vector(23 downto 0) := X"100000";
	signal hsize : unsigned(11 downto 0) := TO_UNSIGNED(640,12);
	signal htotal : unsigned(11 downto 0) := TO_UNSIGNED(800,12);
	signal hbstart : unsigned(11 downto 0) := TO_UNSIGNED(656,12);
	signal hbstop : unsigned(11 downto 0) := TO_UNSIGNED(752,12);
	signal vsize : unsigned(11 downto 0) := TO_UNSIGNED(480,12);
	signal vtotal : unsigned(11 downto 0) := TO_UNSIGNED(525,12);
	signal vbstart : unsigned(11 downto 0) := TO_UNSIGNED(500,12);
	signal vbstop : unsigned(11 downto 0) := TO_UNSIGNED(502,12);

	signal sprite0_pointer : std_logic_vector(23 downto 0) := X"000000";
	signal sprite0_xpos : unsigned(11 downto 0);
	signal sprite0_ypos : unsigned(11 downto 0);
	signal sprite0_data : std_logic_vector(3 downto 0);
	signal set_sprite0 : std_logic;
	signal sprite0_req : std_logic;
	
	signal currentX : unsigned(11 downto 0);
	signal currentY : unsigned(11 downto 0);
	signal end_of_pixel : std_logic;
	signal vga_newframe : std_logic;
	signal vgacache_req : std_logic;
	signal vgadata : std_logic_vector(15 downto 0);
	signal oddframe : std_logic;	-- Toggled each frame, used for dithering

	signal ored : unsigned(5 downto 0);
	signal ogreen : unsigned(5 downto 0);
	signal oblue : unsigned(5 downto 0);
	signal dither : unsigned(5 downto 0);
	signal sprite_col : unsigned(3 downto 0);

	signal chargen_addr : std_logic_vector(10 downto 0);
	signal chargen_datain : std_logic_vector(7 downto 0);
	signal chargen_dataout : std_logic_vector(7 downto 0);
	signal chargen_window : std_logic := '0';
	signal chargen_pixel : std_logic := '0';
	signal chargen_rw : std_logic :='1';

	type charramstates is (writeupperbyte,readupperbyte1,readupperbyte2,writelowerbyte,readlowerbyte1,readlowerbyte2);
	signal charramstate : charramstates;			

begin

	red <= ored(5 downto 2);
	green <= ogreen(5 downto 2);
	blue <= oblue(5 downto 2);

	myVgaMaster : entity work.video_vga_master
		generic map (
			clkDivBits => 4
		)
		port map (
			clk => clk,
			clkDiv => X"3",	-- 100 Mhz / (3+1) = 25 Mhz
--			clkDiv => X"4",	-- 125 Mhz / (4+1) = 25 Mhz

			hSync => hsync,
			vSync => vsync,

			endOfPixel => end_of_pixel,
			endOfLine => open,
			endOfFrame => open,
			currentX => currentX,
			currentY => currentY,

			-- Setup 640x480@60hz needs ~25 Mhz
			hSyncPol => '0',
			vSyncPol => '0',
			xSize => htotal,
			ySize => vtotal,
			xSyncFr => hbstart,
			xSyncTo => hbstop,
			ySyncFr => vbstart, -- Sync pulse 2
			ySyncTo => vbstop
		);		

	myvgacache : entity work.vgacache
		port map(
			clk => clk,
			reset => reset,

			addrin => vga_pointer,
--			idle => sdr_reservebank,

			vga_req => vgacache_req,
			data_out => vgadata,
			setvga => vga_newframe,

			sprite0_out => sprite0_data,
			setsprite0 => set_sprite0,
			sprite0_req => sprite0_req,

			addrout => sdr_addrout,
			data_in => sdr_datain,
			fill => sdr_fill,
			req => sdr_req,
--			reservebank => sdr_reservebank,
--			reservebank => open,
			reserveaddr => sdr_reserveaddr
		);

	mychargen : entity work.charactergenerator
		generic map (
			xstart => 16,
			xstop => 624,
			ystart => 256,
			ystop => 464,
			border => 7
		)
		port map (
			clk => clk,
			reset => reset,
			xpos => currentX(9 downto 0),
			ypos => currentY(9 downto 0),
			pixel_clock => end_of_pixel,
			pixel => chargen_pixel,
			window => chargen_window,
			-- Char RAM access.
			addrin => chargen_addr,
			datain => chargen_datain,
			dataout => chargen_dataout,
			rw => chargen_rw
		);

	-- Handle CPU access to hardware registers
	
	process(clk,reset)
	begin
		if reset='0' then
			htotal <= TO_UNSIGNED(800,12);
			vtotal <= TO_UNSIGNED(525,12);
			hbstart <= TO_UNSIGNED(656,12);
			hbstop <= TO_UNSIGNED(752,12);
			vbstart <= TO_UNSIGNED(500,12);
			vbstop <= TO_UNSIGNED(502,12);
			reg_data_out<=X"0000";
			sprite0_xpos<=X"000";
			sprite0_ypos<=X"000";
			chargen_addr<="00000000000";
		elsif rising_edge(clk) then
			reg_dtack<='1';
			chargen_rw<='1';

			charramstate<=writeupperbyte; -- Reset state machine.
			if reg_addr_in(11)='1' then	-- Character RAM access
				-- Need to deal with both word and byte reads/writes.
				-- We do one read and one write to both bytes on a 4-step cycle.
				case charramstate is
					when writeupperbyte =>
						if reg_req='1' then
							chargen_addr<=reg_addr_in(10 downto 1) & '0';	-- Upper byte
							chargen_datain<=reg_data_in(15 downto 8);
							if reg_rw='0' and reg_uds='0' then
								chargen_rw<='0';
							end if;
							charramstate<=readupperbyte1;
						end if;
					when readupperbyte1 =>
						charramstate<=readupperbyte2;	-- delay for data
					when readupperbyte2 =>			
						reg_data_out(15 downto 8)<=chargen_dataout;
						charramstate<=writelowerbyte;
					when writelowerbyte =>
						chargen_addr<=reg_addr_in(10 downto 1) & '1';	-- lower byte
						chargen_datain<=reg_data_in(7 downto 0);
						if reg_rw='0' and reg_lds='0' then
							chargen_rw<='0';
						end if;
						charramstate<=readlowerbyte1;
					when readlowerbyte1 =>
						charramstate<=readlowerbyte2;	-- delay for data
					when readlowerbyte2 =>
						reg_data_out(7 downto 0)<=chargen_dataout;
						reg_dtack<='0';
				end case;
			elsif reg_req='1' then
				case reg_addr_in is
					when X"000" =>
	--					reg_data_out<=X"00"&framebuffer_pointer(23 downto 16);
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							framebuffer_pointer(23 downto 16) <= reg_data_in(7 downto 0);
						end if;
					when X"002" =>
	--					reg_data_out<=framebuffer_pointer(15 downto 0);
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							framebuffer_pointer(15 downto 0) <= reg_data_in;
						end if;
					when X"100" =>
	--					reg_data_out<=X"00"&sprite0_pointer(23 downto 16);
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							sprite0_pointer(23 downto 16) <= reg_data_in(7 downto 0);
						end if;
					when X"102" =>
	--					reg_data_out<=sprite0_pointer(15 downto 0);
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							sprite0_pointer(15 downto 0) <= reg_data_in;
						end if;
					when X"104" =>
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							sprite0_xpos <= unsigned(reg_data_in(11 downto 0));
						end if;
					when X"106" =>
						if reg_rw='0' and reg_uds='0' and reg_lds='0' then
							sprite0_ypos <= unsigned(reg_data_in(11 downto 0));
						end if;
					when others =>
						reg_data_out<=X"0000";
				end case;
				reg_dtack<='0';
			end if;
-- FBPTH equ $0000	; Framebuffer pointer - must be 64-bit aligned.
-- FBPTL equ $0002

--     4   Even row modulo
--     6   Odd row modulo (allows scandoubling)

--     8  HTotal
--     A  HSize (typically 640)
--     C  HBStart
--     E  HBStop

--    10  VTotal
--    12  VSize (typically 480)
--    14  VBStart
--    16  VBStop

--    18  Control:
--     0  Visible
--     1  Resolution - high, low  - alternatively could make pixel clock programmable...
--     7  Character overlay on/off

-- SP0PTH equ $0100 ; Pointer to sprite 0's data - must be 64-bit aligned.
-- SP0PTL equ $0102
-- SP0XPOS	equ $0104
-- SP0YPOS equ $0106


		end if;
	end process;

	
	-- Sprite positions
	process(clk, reset, currentX, currentY)
	begin
		if rising_edge(clk) then
			sprite0_req<='0';
			if currentX>=sprite0_xpos and currentX-sprite0_xpos<16
						and currentY>=sprite0_ypos and currentY-sprite0_ypos<16 then	
				if end_of_pixel='1' then
					sprite_col<=unsigned(sprite0_data);
					sprite0_req<='1';
				end if;
			else
				sprite_col<="0000";
			end if;
		end if;
	end process;
	
	
	process(clk, reset,currentX, currentY)
	begin
		if rising_edge(clk) then
			sdr_refresh <='0';
			if end_of_pixel='1' and currentX=hsize then
				sdr_refresh<='1';
			end if;
		end if;
		
		if reset='0' then
			vgacache_req <='0';
			sdr_reservebank<='1';
		elsif rising_edge(clk) then
			vblank_int<='0';
			vgacache_req<='0';
			vga_newframe<='0';
			vgacache_req<='0';
			set_sprite0<='0';
			if end_of_pixel='1' then
				sdr_reservebank<='1';
			-- Dither: bit 1: temporal dithering, alternate lines swapped each frame
				--         bit 0: spatial dithering, alternate pixels
				dither<="0000" & (currentY(0) xor oddframe) & (currentX(0) xor currentY(0));

				if currentX<640 and currentY<480 then
					-- Request next pixel from VGA cache
					vgacache_req<='1';

					-- Now dither the pixel.  If we're drawing a pixel from the character
					-- generator or sprites, or the pixel is already at max, we don't dither. (Avoids overflow)
					if sprite_col(3)='1' then
						ored <= sprite_col(2) & sprite_col(2) & sprite_col(2) & 
							sprite_col(2) & sprite_col(2) & sprite_col(2);
					elsif chargen_pixel='1' or (chargen_window='0' and vgadata(15 downto 12)="1111") then
						ored <= "111111";
					elsif chargen_window='1' then
						ored <= unsigned('0'&vgadata(15 downto 11)) + dither;
					else
						ored <= unsigned(vgadata(15 downto 11)&'0') + dither;
					end if;

					if sprite_col(3)='1' then
						ogreen <= sprite_col(1) & sprite_col(1) & sprite_col(1) & 
							sprite_col(1) & sprite_col(1) & sprite_col(1);
					elsif chargen_pixel='1' or (chargen_window='0' and vgadata(10 downto 7)="1111") then
						ogreen <= "111111";
					elsif chargen_window='1' then
						ogreen <= unsigned('0'&vgadata(10 downto 6)) + dither;
					else
						ogreen <= unsigned(vgadata(10 downto 5)) + dither;
					end if;

					if sprite_col(3)='1' then
						oblue <= sprite_col(0) & sprite_col(0) & sprite_col(0) & 
							sprite_col(0) & sprite_col(0) & sprite_col(0);
					elsif chargen_pixel='1' or (chargen_window='0' and vgadata(4 downto 1)="1111") then
						oblue <= "111111";
					elsif chargen_window='1' then
						oblue <= unsigned('0'&vgadata(4 downto 0)) + dither;
					else
						oblue <= unsigned(vgadata(4 downto 0)&'0') + dither;
					end if;

				else
					ored<="000000"; -- need to set black during sync periods.
					ogreen<="000000";
					oblue<="000000";
					if currentY=vsize and currentX=0 then
						oddframe<=not oddframe;
						vga_pointer<=framebuffer_pointer;
						vga_newframe<='1';
						vblank_int<='1';
					end if;

					if currentY=vtotal and currentX=0 then
						vga_pointer<=sprite0_pointer;
						set_sprite0<='1';
					end if;
					
--					if currentX>(hsize+12) and currentX<(htotal - 4) then	-- Signal to SDRAM controller that we're
					if currentX<(htotal - 6) then	-- Signal to SDRAM controller that we're
						sdr_reservebank<='0'; -- in blank areas, so there's no need to keep slot 2 off the next bank.
					end if;
				end if;
			end if;
		end if;
	end process;
		
end architecture;
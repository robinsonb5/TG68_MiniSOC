library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"33",
    49 => x"fc",
    50 => x"00",
    51 => x"01",
    52 => x"81",
    53 => x"00",
    54 => x"00",
    55 => x"04",
    56 => x"41",
    57 => x"fa",
    58 => x"00",
    59 => x"80",
    60 => x"61",
    61 => x"00",
    62 => x"02",
    63 => x"e4",
    64 => x"33",
    65 => x"fc",
    66 => x"0f",
    67 => x"00",
    68 => x"81",
    69 => x"00",
    70 => x"00",
    71 => x"06",
    72 => x"2e",
    73 => x"3c",
    74 => x"00",
    75 => x"00",
    76 => x"07",
    77 => x"ff",
    78 => x"41",
    79 => x"f9",
    80 => x"80",
    81 => x"00",
    82 => x"08",
    83 => x"00",
    84 => x"10",
    85 => x"fc",
    86 => x"00",
    87 => x"20",
    88 => x"51",
    89 => x"cf",
    90 => x"ff",
    91 => x"fa",
    92 => x"23",
    93 => x"fc",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"7f",
   100 => x"00",
   101 => x"52",
   102 => x"41",
   103 => x"fa",
   104 => x"00",
   105 => x"52",
   106 => x"61",
   107 => x"00",
   108 => x"06",
   109 => x"c6",
   110 => x"61",
   111 => x"00",
   112 => x"0a",
   113 => x"f8",
   114 => x"4a",
   115 => x"80",
   116 => x"67",
   117 => x"0a",
   118 => x"41",
   119 => x"fa",
   120 => x"00",
   121 => x"76",
   122 => x"61",
   123 => x"00",
   124 => x"06",
   125 => x"b6",
   126 => x"60",
   127 => x"fe",
   128 => x"41",
   129 => x"fa",
   130 => x"00",
   131 => x"55",
   132 => x"61",
   133 => x"00",
   134 => x"06",
   135 => x"ac",
   136 => x"61",
   137 => x"00",
   138 => x"02",
   139 => x"b8",
   140 => x"4b",
   141 => x"f9",
   142 => x"80",
   143 => x"00",
   144 => x"08",
   145 => x"00",
   146 => x"33",
   147 => x"fc",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"7f",
   152 => x"00",
   153 => x"0c",
   154 => x"30",
   155 => x"39",
   156 => x"81",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"08",
   161 => x"00",
   162 => x"00",
   163 => x"09",
   164 => x"67",
   165 => x"f4",
   166 => x"1a",
   167 => x"c0",
   168 => x"22",
   169 => x"0d",
   170 => x"82",
   171 => x"b8",
   172 => x"08",
   173 => x"00",
   174 => x"c2",
   175 => x"b8",
   176 => x"ef",
   177 => x"ff",
   178 => x"2a",
   179 => x"41",
   180 => x"61",
   181 => x"00",
   182 => x"00",
   183 => x"80",
   184 => x"60",
   185 => x"e0",
   186 => x"43",
   187 => x"6f",
   188 => x"6e",
   189 => x"64",
   190 => x"75",
   191 => x"63",
   192 => x"74",
   193 => x"69",
   194 => x"6e",
   195 => x"67",
   196 => x"20",
   197 => x"73",
   198 => x"61",
   199 => x"6e",
   200 => x"69",
   201 => x"74",
   202 => x"79",
   203 => x"20",
   204 => x"63",
   205 => x"68",
   206 => x"65",
   207 => x"63",
   208 => x"6b",
   209 => x"2e",
   210 => x"2e",
   211 => x"2e",
   212 => x"0d",
   213 => x"0a",
   214 => x"00",
   215 => x"53",
   216 => x"61",
   217 => x"6e",
   218 => x"69",
   219 => x"74",
   220 => x"79",
   221 => x"20",
   222 => x"63",
   223 => x"68",
   224 => x"65",
   225 => x"63",
   226 => x"6b",
   227 => x"20",
   228 => x"70",
   229 => x"61",
   230 => x"73",
   231 => x"73",
   232 => x"65",
   233 => x"64",
   234 => x"2e",
   235 => x"0d",
   236 => x"0a",
   237 => x"00",
   238 => x"53",
   239 => x"61",
   240 => x"6e",
   241 => x"69",
   242 => x"74",
   243 => x"79",
   244 => x"20",
   245 => x"63",
   246 => x"68",
   247 => x"65",
   248 => x"63",
   249 => x"6b",
   250 => x"20",
   251 => x"66",
   252 => x"61",
   253 => x"69",
   254 => x"6c",
   255 => x"65",
   256 => x"64",
   257 => x"2e",
   258 => x"0d",
   259 => x"0a",
   260 => x"00",
   261 => x"00",
   262 => x"c0",
   263 => x"bc",
   264 => x"00",
   265 => x"00",
   266 => x"00",
   267 => x"df",
   268 => x"90",
   269 => x"3c",
   270 => x"00",
   271 => x"37",
   272 => x"6a",
   273 => x"04",
   274 => x"d0",
   275 => x"3c",
   276 => x"00",
   277 => x"27",
   278 => x"e9",
   279 => x"8e",
   280 => x"8c",
   281 => x"00",
   282 => x"20",
   283 => x"86",
   284 => x"4e",
   285 => x"75",
   286 => x"c0",
   287 => x"bc",
   288 => x"00",
   289 => x"00",
   290 => x"00",
   291 => x"df",
   292 => x"90",
   293 => x"3c",
   294 => x"00",
   295 => x"37",
   296 => x"6a",
   297 => x"04",
   298 => x"d0",
   299 => x"3c",
   300 => x"00",
   301 => x"27",
   302 => x"e9",
   303 => x"0f",
   304 => x"8e",
   305 => x"00",
   306 => x"10",
   307 => x"87",
   308 => x"4e",
   309 => x"75",
   310 => x"52",
   311 => x"79",
   312 => x"00",
   313 => x"7f",
   314 => x"00",
   315 => x"0c",
   316 => x"b0",
   317 => x"3c",
   318 => x"00",
   319 => x"53",
   320 => x"66",
   321 => x"2a",
   322 => x"33",
   323 => x"fc",
   324 => x"ff",
   325 => x"ff",
   326 => x"81",
   327 => x"00",
   328 => x"00",
   329 => x"06",
   330 => x"72",
   331 => x"00",
   332 => x"2e",
   333 => x"01",
   334 => x"2c",
   335 => x"01",
   336 => x"33",
   337 => x"c1",
   338 => x"00",
   339 => x"7f",
   340 => x"00",
   341 => x"0c",
   342 => x"23",
   343 => x"c1",
   344 => x"00",
   345 => x"7f",
   346 => x"00",
   347 => x"08",
   348 => x"23",
   349 => x"c1",
   350 => x"00",
   351 => x"7f",
   352 => x"00",
   353 => x"04",
   354 => x"23",
   355 => x"c1",
   356 => x"00",
   357 => x"7f",
   358 => x"00",
   359 => x"10",
   360 => x"60",
   361 => x"00",
   362 => x"01",
   363 => x"72",
   364 => x"2c",
   365 => x"39",
   366 => x"00",
   367 => x"7f",
   368 => x"00",
   369 => x"20",
   370 => x"2e",
   371 => x"39",
   372 => x"00",
   373 => x"7f",
   374 => x"00",
   375 => x"1c",
   376 => x"0c",
   377 => x"79",
   378 => x"00",
   379 => x"01",
   380 => x"00",
   381 => x"7f",
   382 => x"00",
   383 => x"0c",
   384 => x"66",
   385 => x"34",
   386 => x"33",
   387 => x"fc",
   388 => x"f0",
   389 => x"00",
   390 => x"81",
   391 => x"00",
   392 => x"00",
   393 => x"06",
   394 => x"41",
   395 => x"f9",
   396 => x"00",
   397 => x"7f",
   398 => x"00",
   399 => x"13",
   400 => x"61",
   401 => x"8c",
   402 => x"22",
   403 => x"39",
   404 => x"00",
   405 => x"7f",
   406 => x"00",
   407 => x"10",
   408 => x"b2",
   409 => x"bc",
   410 => x"00",
   411 => x"00",
   412 => x"00",
   413 => x"03",
   414 => x"6f",
   415 => x"08",
   416 => x"72",
   417 => x"0a",
   418 => x"92",
   419 => x"b9",
   420 => x"00",
   421 => x"7f",
   422 => x"00",
   423 => x"10",
   424 => x"52",
   425 => x"81",
   426 => x"e3",
   427 => x"89",
   428 => x"23",
   429 => x"c1",
   430 => x"00",
   431 => x"7f",
   432 => x"00",
   433 => x"14",
   434 => x"60",
   435 => x"00",
   436 => x"01",
   437 => x"28",
   438 => x"33",
   439 => x"f9",
   440 => x"00",
   441 => x"7f",
   442 => x"00",
   443 => x"12",
   444 => x"81",
   445 => x"00",
   446 => x"00",
   447 => x"06",
   448 => x"4a",
   449 => x"b9",
   450 => x"00",
   451 => x"7f",
   452 => x"00",
   453 => x"10",
   454 => x"67",
   455 => x"00",
   456 => x"01",
   457 => x"14",
   458 => x"0c",
   459 => x"b9",
   460 => x"00",
   461 => x"00",
   462 => x"00",
   463 => x"09",
   464 => x"00",
   465 => x"7f",
   466 => x"00",
   467 => x"10",
   468 => x"6e",
   469 => x"00",
   470 => x"00",
   471 => x"c0",
   472 => x"0c",
   473 => x"79",
   474 => x"00",
   475 => x"03",
   476 => x"00",
   477 => x"7f",
   478 => x"00",
   479 => x"0c",
   480 => x"6e",
   481 => x"16",
   482 => x"33",
   483 => x"fc",
   484 => x"0f",
   485 => x"00",
   486 => x"81",
   487 => x"00",
   488 => x"00",
   489 => x"06",
   490 => x"41",
   491 => x"f9",
   492 => x"00",
   493 => x"7f",
   494 => x"00",
   495 => x"07",
   496 => x"61",
   497 => x"00",
   498 => x"ff",
   499 => x"2c",
   500 => x"60",
   501 => x"00",
   502 => x"00",
   503 => x"e6",
   504 => x"22",
   505 => x"39",
   506 => x"00",
   507 => x"7f",
   508 => x"00",
   509 => x"14",
   510 => x"56",
   511 => x"41",
   512 => x"34",
   513 => x"39",
   514 => x"00",
   515 => x"7f",
   516 => x"00",
   517 => x"0c",
   518 => x"b4",
   519 => x"41",
   520 => x"6e",
   521 => x"20",
   522 => x"41",
   523 => x"f9",
   524 => x"00",
   525 => x"7f",
   526 => x"00",
   527 => x"08",
   528 => x"61",
   529 => x"00",
   530 => x"fe",
   531 => x"f4",
   532 => x"33",
   533 => x"f9",
   534 => x"00",
   535 => x"7f",
   536 => x"00",
   537 => x"0a",
   538 => x"81",
   539 => x"00",
   540 => x"00",
   541 => x"06",
   542 => x"33",
   543 => x"fc",
   544 => x"00",
   545 => x"01",
   546 => x"00",
   547 => x"7f",
   548 => x"00",
   549 => x"18",
   550 => x"60",
   551 => x"00",
   552 => x"00",
   553 => x"b4",
   554 => x"0c",
   555 => x"b9",
   556 => x"00",
   557 => x"00",
   558 => x"00",
   559 => x"03",
   560 => x"00",
   561 => x"7f",
   562 => x"00",
   563 => x"10",
   564 => x"6e",
   565 => x"60",
   566 => x"33",
   567 => x"fc",
   568 => x"00",
   569 => x"0f",
   570 => x"81",
   571 => x"00",
   572 => x"00",
   573 => x"06",
   574 => x"22",
   575 => x"39",
   576 => x"00",
   577 => x"7f",
   578 => x"00",
   579 => x"04",
   580 => x"e3",
   581 => x"89",
   582 => x"52",
   583 => x"81",
   584 => x"34",
   585 => x"39",
   586 => x"00",
   587 => x"7f",
   588 => x"00",
   589 => x"0c",
   590 => x"b4",
   591 => x"41",
   592 => x"6e",
   593 => x"2a",
   594 => x"20",
   595 => x"79",
   596 => x"00",
   597 => x"7f",
   598 => x"00",
   599 => x"08",
   600 => x"61",
   601 => x"00",
   602 => x"fe",
   603 => x"c4",
   604 => x"32",
   605 => x"39",
   606 => x"00",
   607 => x"7f",
   608 => x"00",
   609 => x"18",
   610 => x"53",
   611 => x"79",
   612 => x"00",
   613 => x"7f",
   614 => x"00",
   615 => x"18",
   616 => x"53",
   617 => x"41",
   618 => x"6a",
   619 => x"70",
   620 => x"52",
   621 => x"b9",
   622 => x"00",
   623 => x"7f",
   624 => x"00",
   625 => x"08",
   626 => x"33",
   627 => x"fc",
   628 => x"00",
   629 => x"01",
   630 => x"00",
   631 => x"7f",
   632 => x"00",
   633 => x"18",
   634 => x"60",
   635 => x"60",
   636 => x"30",
   637 => x"39",
   638 => x"00",
   639 => x"7f",
   640 => x"00",
   641 => x"18",
   642 => x"52",
   643 => x"40",
   644 => x"c0",
   645 => x"7c",
   646 => x"00",
   647 => x"01",
   648 => x"67",
   649 => x"52",
   650 => x"20",
   651 => x"79",
   652 => x"00",
   653 => x"7f",
   654 => x"00",
   655 => x"08",
   656 => x"e5",
   657 => x"88",
   658 => x"e1",
   659 => x"2f",
   660 => x"10",
   661 => x"87",
   662 => x"33",
   663 => x"fc",
   664 => x"f0",
   665 => x"f0",
   666 => x"81",
   667 => x"00",
   668 => x"00",
   669 => x"06",
   670 => x"0c",
   671 => x"b9",
   672 => x"00",
   673 => x"00",
   674 => x"00",
   675 => x"07",
   676 => x"00",
   677 => x"7f",
   678 => x"00",
   679 => x"10",
   680 => x"6d",
   681 => x"32",
   682 => x"33",
   683 => x"fc",
   684 => x"f0",
   685 => x"0f",
   686 => x"81",
   687 => x"00",
   688 => x"00",
   689 => x"06",
   690 => x"0c",
   691 => x"b9",
   692 => x"00",
   693 => x"00",
   694 => x"00",
   695 => x"09",
   696 => x"00",
   697 => x"7f",
   698 => x"00",
   699 => x"10",
   700 => x"6e",
   701 => x"1e",
   702 => x"33",
   703 => x"fc",
   704 => x"ff",
   705 => x"f0",
   706 => x"81",
   707 => x"00",
   708 => x"00",
   709 => x"06",
   710 => x"41",
   711 => x"fa",
   712 => x"00",
   713 => x"22",
   714 => x"61",
   715 => x"56",
   716 => x"2e",
   717 => x"b9",
   718 => x"00",
   719 => x"7f",
   720 => x"00",
   721 => x"08",
   722 => x"08",
   723 => x"b9",
   724 => x"00",
   725 => x"00",
   726 => x"81",
   727 => x"00",
   728 => x"00",
   729 => x"04",
   730 => x"4e",
   731 => x"75",
   732 => x"23",
   733 => x"c6",
   734 => x"00",
   735 => x"7f",
   736 => x"00",
   737 => x"20",
   738 => x"23",
   739 => x"c7",
   740 => x"00",
   741 => x"7f",
   742 => x"00",
   743 => x"1c",
   744 => x"4e",
   745 => x"75",
   746 => x"46",
   747 => x"69",
   748 => x"72",
   749 => x"6d",
   750 => x"77",
   751 => x"61",
   752 => x"72",
   753 => x"65",
   754 => x"20",
   755 => x"72",
   756 => x"65",
   757 => x"63",
   758 => x"65",
   759 => x"69",
   760 => x"76",
   761 => x"65",
   762 => x"64",
   763 => x"20",
   764 => x"2d",
   765 => x"20",
   766 => x"6c",
   767 => x"61",
   768 => x"75",
   769 => x"6e",
   770 => x"63",
   771 => x"68",
   772 => x"69",
   773 => x"6e",
   774 => x"67",
   775 => x"0d",
   776 => x"0a",
   777 => x"00",
   778 => x"48",
   779 => x"40",
   780 => x"30",
   781 => x"39",
   782 => x"81",
   783 => x"00",
   784 => x"00",
   785 => x"00",
   786 => x"08",
   787 => x"00",
   788 => x"00",
   789 => x"08",
   790 => x"67",
   791 => x"f4",
   792 => x"48",
   793 => x"40",
   794 => x"33",
   795 => x"c0",
   796 => x"81",
   797 => x"00",
   798 => x"00",
   799 => x"00",
   800 => x"4e",
   801 => x"75",
   802 => x"2f",
   803 => x"00",
   804 => x"70",
   805 => x"00",
   806 => x"30",
   807 => x"39",
   808 => x"81",
   809 => x"00",
   810 => x"00",
   811 => x"00",
   812 => x"08",
   813 => x"00",
   814 => x"00",
   815 => x"08",
   816 => x"67",
   817 => x"f4",
   818 => x"10",
   819 => x"18",
   820 => x"67",
   821 => x"08",
   822 => x"33",
   823 => x"c0",
   824 => x"81",
   825 => x"00",
   826 => x"00",
   827 => x"00",
   828 => x"60",
   829 => x"e8",
   830 => x"20",
   831 => x"1f",
   832 => x"4e",
   833 => x"75",
   834 => x"33",
   835 => x"fc",
   836 => x"00",
   837 => x"01",
   838 => x"81",
   839 => x"00",
   840 => x"00",
   841 => x"06",
   842 => x"41",
   843 => x"fa",
   844 => x"01",
   845 => x"fa",
   846 => x"61",
   847 => x"00",
   848 => x"03",
   849 => x"e2",
   850 => x"61",
   851 => x"00",
   852 => x"02",
   853 => x"60",
   854 => x"66",
   855 => x"5c",
   856 => x"33",
   857 => x"fc",
   858 => x"00",
   859 => x"02",
   860 => x"81",
   861 => x"00",
   862 => x"00",
   863 => x"06",
   864 => x"33",
   865 => x"fc",
   866 => x"00",
   867 => x"40",
   868 => x"00",
   869 => x"7f",
   870 => x"00",
   871 => x"26",
   872 => x"61",
   873 => x"00",
   874 => x"04",
   875 => x"8a",
   876 => x"67",
   877 => x"0c",
   878 => x"42",
   879 => x"79",
   880 => x"00",
   881 => x"7f",
   882 => x"00",
   883 => x"26",
   884 => x"61",
   885 => x"00",
   886 => x"04",
   887 => x"7e",
   888 => x"66",
   889 => x"28",
   890 => x"33",
   891 => x"fc",
   892 => x"00",
   893 => x"03",
   894 => x"81",
   895 => x"00",
   896 => x"00",
   897 => x"06",
   898 => x"61",
   899 => x"00",
   900 => x"05",
   901 => x"f8",
   902 => x"43",
   903 => x"fa",
   904 => x"00",
   905 => x"57",
   906 => x"61",
   907 => x"00",
   908 => x"06",
   909 => x"48",
   910 => x"67",
   911 => x"12",
   912 => x"41",
   913 => x"fa",
   914 => x"00",
   915 => x"47",
   916 => x"61",
   917 => x"00",
   918 => x"03",
   919 => x"9c",
   920 => x"30",
   921 => x"7c",
   922 => x"20",
   923 => x"00",
   924 => x"61",
   925 => x"00",
   926 => x"04",
   927 => x"02",
   928 => x"4e",
   929 => x"75",
   930 => x"33",
   931 => x"fc",
   932 => x"f0",
   933 => x"03",
   934 => x"81",
   935 => x"00",
   936 => x"00",
   937 => x"06",
   938 => x"41",
   939 => x"fa",
   940 => x"00",
   941 => x"29",
   942 => x"61",
   943 => x"00",
   944 => x"03",
   945 => x"82",
   946 => x"4e",
   947 => x"75",
   948 => x"33",
   949 => x"fc",
   950 => x"f0",
   951 => x"02",
   952 => x"81",
   953 => x"00",
   954 => x"00",
   955 => x"06",
   956 => x"41",
   957 => x"fa",
   958 => x"00",
   959 => x"08",
   960 => x"61",
   961 => x"00",
   962 => x"03",
   963 => x"70",
   964 => x"4e",
   965 => x"75",
   966 => x"53",
   967 => x"44",
   968 => x"20",
   969 => x"69",
   970 => x"6e",
   971 => x"69",
   972 => x"74",
   973 => x"20",
   974 => x"66",
   975 => x"61",
   976 => x"69",
   977 => x"6c",
   978 => x"65",
   979 => x"64",
   980 => x"00",
   981 => x"6e",
   982 => x"6f",
   983 => x"74",
   984 => x"20",
   985 => x"66",
   986 => x"6f",
   987 => x"75",
   988 => x"6e",
   989 => x"64",
   990 => x"20",
   991 => x"42",
   992 => x"4f",
   993 => x"4f",
   994 => x"54",
   995 => x"20",
   996 => x"20",
   997 => x"20",
   998 => x"20",
   999 => x"53",
  1000 => x"52",
  1001 => x"45",
  1002 => x"00",
  1003 => x"00",
  1004 => x"33",
  1005 => x"fc",
  1006 => x"01",
  1007 => x"00",
  1008 => x"81",
  1009 => x"00",
  1010 => x"00",
  1011 => x"06",
  1012 => x"41",
  1013 => x"f9",
  1014 => x"00",
  1015 => x"7f",
  1016 => x"00",
  1017 => x"56",
  1018 => x"61",
  1019 => x"00",
  1020 => x"00",
  1021 => x"c4",
  1022 => x"66",
  1023 => x"68",
  1024 => x"33",
  1025 => x"fc",
  1026 => x"01",
  1027 => x"01",
  1028 => x"81",
  1029 => x"00",
  1030 => x"00",
  1031 => x"06",
  1032 => x"32",
  1033 => x"3c",
  1034 => x"4e",
  1035 => x"20",
  1036 => x"53",
  1037 => x"41",
  1038 => x"67",
  1039 => x"44",
  1040 => x"33",
  1041 => x"fc",
  1042 => x"01",
  1043 => x"02",
  1044 => x"81",
  1045 => x"00",
  1046 => x"00",
  1047 => x"06",
  1048 => x"33",
  1049 => x"7c",
  1050 => x"00",
  1051 => x"ff",
  1052 => x"00",
  1053 => x"24",
  1054 => x"30",
  1055 => x"29",
  1056 => x"00",
  1057 => x"24",
  1058 => x"b0",
  1059 => x"3c",
  1060 => x"00",
  1061 => x"fe",
  1062 => x"66",
  1063 => x"e4",
  1064 => x"30",
  1065 => x"29",
  1066 => x"01",
  1067 => x"00",
  1068 => x"32",
  1069 => x"3c",
  1070 => x"00",
  1071 => x"7f",
  1072 => x"20",
  1073 => x"29",
  1074 => x"01",
  1075 => x"00",
  1076 => x"20",
  1077 => x"c0",
  1078 => x"51",
  1079 => x"c9",
  1080 => x"ff",
  1081 => x"f8",
  1082 => x"30",
  1083 => x"29",
  1084 => x"00",
  1085 => x"24",
  1086 => x"33",
  1087 => x"7c",
  1088 => x"00",
  1089 => x"00",
  1090 => x"00",
  1091 => x"22",
  1092 => x"33",
  1093 => x"fc",
  1094 => x"01",
  1095 => x"03",
  1096 => x"81",
  1097 => x"00",
  1098 => x"00",
  1099 => x"06",
  1100 => x"41",
  1101 => x"e8",
  1102 => x"fe",
  1103 => x"00",
  1104 => x"70",
  1105 => x"00",
  1106 => x"4e",
  1107 => x"75",
  1108 => x"33",
  1109 => x"fc",
  1110 => x"f1",
  1111 => x"02",
  1112 => x"81",
  1113 => x"00",
  1114 => x"00",
  1115 => x"06",
  1116 => x"41",
  1117 => x"fa",
  1118 => x"01",
  1119 => x"38",
  1120 => x"61",
  1121 => x"00",
  1122 => x"02",
  1123 => x"d0",
  1124 => x"70",
  1125 => x"fe",
  1126 => x"4e",
  1127 => x"75",
  1128 => x"33",
  1129 => x"fc",
  1130 => x"f1",
  1131 => x"03",
  1132 => x"81",
  1133 => x"00",
  1134 => x"00",
  1135 => x"06",
  1136 => x"41",
  1137 => x"fa",
  1138 => x"01",
  1139 => x"0c",
  1140 => x"61",
  1141 => x"00",
  1142 => x"02",
  1143 => x"bc",
  1144 => x"70",
  1145 => x"ff",
  1146 => x"4e",
  1147 => x"75",
  1148 => x"22",
  1149 => x"3c",
  1150 => x"00",
  1151 => x"95",
  1152 => x"00",
  1153 => x"40",
  1154 => x"70",
  1155 => x"00",
  1156 => x"60",
  1157 => x"40",
  1158 => x"22",
  1159 => x"3c",
  1160 => x"00",
  1161 => x"ff",
  1162 => x"00",
  1163 => x"41",
  1164 => x"70",
  1165 => x"00",
  1166 => x"60",
  1167 => x"36",
  1168 => x"22",
  1169 => x"3c",
  1170 => x"00",
  1171 => x"87",
  1172 => x"00",
  1173 => x"48",
  1174 => x"20",
  1175 => x"3c",
  1176 => x"00",
  1177 => x"00",
  1178 => x"01",
  1179 => x"aa",
  1180 => x"60",
  1181 => x"28",
  1182 => x"22",
  1183 => x"3c",
  1184 => x"00",
  1185 => x"87",
  1186 => x"00",
  1187 => x"69",
  1188 => x"20",
  1189 => x"3c",
  1190 => x"40",
  1191 => x"00",
  1192 => x"00",
  1193 => x"00",
  1194 => x"60",
  1195 => x"1a",
  1196 => x"22",
  1197 => x"3c",
  1198 => x"00",
  1199 => x"ff",
  1200 => x"00",
  1201 => x"77",
  1202 => x"70",
  1203 => x"00",
  1204 => x"60",
  1205 => x"10",
  1206 => x"22",
  1207 => x"3c",
  1208 => x"00",
  1209 => x"ff",
  1210 => x"00",
  1211 => x"7a",
  1212 => x"70",
  1213 => x"00",
  1214 => x"60",
  1215 => x"06",
  1216 => x"22",
  1217 => x"3c",
  1218 => x"00",
  1219 => x"ff",
  1220 => x"00",
  1221 => x"51",
  1222 => x"43",
  1223 => x"f9",
  1224 => x"81",
  1225 => x"00",
  1226 => x"00",
  1227 => x"00",
  1228 => x"33",
  1229 => x"7c",
  1230 => x"00",
  1231 => x"ff",
  1232 => x"00",
  1233 => x"24",
  1234 => x"3f",
  1235 => x"69",
  1236 => x"00",
  1237 => x"24",
  1238 => x"ff",
  1239 => x"fe",
  1240 => x"33",
  1241 => x"7c",
  1242 => x"00",
  1243 => x"01",
  1244 => x"00",
  1245 => x"22",
  1246 => x"33",
  1247 => x"7c",
  1248 => x"00",
  1249 => x"ff",
  1250 => x"00",
  1251 => x"24",
  1252 => x"33",
  1253 => x"41",
  1254 => x"00",
  1255 => x"24",
  1256 => x"48",
  1257 => x"41",
  1258 => x"4a",
  1259 => x"79",
  1260 => x"00",
  1261 => x"7f",
  1262 => x"00",
  1263 => x"24",
  1264 => x"67",
  1265 => x"16",
  1266 => x"e1",
  1267 => x"98",
  1268 => x"33",
  1269 => x"40",
  1270 => x"00",
  1271 => x"24",
  1272 => x"e1",
  1273 => x"98",
  1274 => x"33",
  1275 => x"40",
  1276 => x"00",
  1277 => x"24",
  1278 => x"e1",
  1279 => x"98",
  1280 => x"33",
  1281 => x"40",
  1282 => x"00",
  1283 => x"24",
  1284 => x"e1",
  1285 => x"98",
  1286 => x"60",
  1287 => x"18",
  1288 => x"d0",
  1289 => x"80",
  1290 => x"48",
  1291 => x"40",
  1292 => x"33",
  1293 => x"40",
  1294 => x"00",
  1295 => x"24",
  1296 => x"48",
  1297 => x"40",
  1298 => x"e1",
  1299 => x"58",
  1300 => x"33",
  1301 => x"40",
  1302 => x"00",
  1303 => x"24",
  1304 => x"e1",
  1305 => x"58",
  1306 => x"33",
  1307 => x"40",
  1308 => x"00",
  1309 => x"24",
  1310 => x"70",
  1311 => x"00",
  1312 => x"33",
  1313 => x"40",
  1314 => x"00",
  1315 => x"24",
  1316 => x"33",
  1317 => x"41",
  1318 => x"00",
  1319 => x"24",
  1320 => x"22",
  1321 => x"3c",
  1322 => x"00",
  1323 => x"00",
  1324 => x"01",
  1325 => x"90",
  1326 => x"53",
  1327 => x"81",
  1328 => x"67",
  1329 => x"10",
  1330 => x"33",
  1331 => x"7c",
  1332 => x"00",
  1333 => x"ff",
  1334 => x"00",
  1335 => x"24",
  1336 => x"30",
  1337 => x"29",
  1338 => x"00",
  1339 => x"24",
  1340 => x"b0",
  1341 => x"3c",
  1342 => x"00",
  1343 => x"ff",
  1344 => x"67",
  1345 => x"ec",
  1346 => x"80",
  1347 => x"00",
  1348 => x"4e",
  1349 => x"75",
  1350 => x"53",
  1351 => x"74",
  1352 => x"61",
  1353 => x"72",
  1354 => x"74",
  1355 => x"20",
  1356 => x"49",
  1357 => x"6e",
  1358 => x"69",
  1359 => x"74",
  1360 => x"0d",
  1361 => x"0a",
  1362 => x"00",
  1363 => x"49",
  1364 => x"6e",
  1365 => x"69",
  1366 => x"74",
  1367 => x"20",
  1368 => x"64",
  1369 => x"6f",
  1370 => x"6e",
  1371 => x"65",
  1372 => x"0d",
  1373 => x"0a",
  1374 => x"00",
  1375 => x"49",
  1376 => x"6e",
  1377 => x"69",
  1378 => x"74",
  1379 => x"20",
  1380 => x"66",
  1381 => x"61",
  1382 => x"69",
  1383 => x"6c",
  1384 => x"75",
  1385 => x"72",
  1386 => x"65",
  1387 => x"0d",
  1388 => x"0a",
  1389 => x"00",
  1390 => x"52",
  1391 => x"65",
  1392 => x"73",
  1393 => x"65",
  1394 => x"74",
  1395 => x"20",
  1396 => x"66",
  1397 => x"61",
  1398 => x"69",
  1399 => x"6c",
  1400 => x"75",
  1401 => x"72",
  1402 => x"65",
  1403 => x"0d",
  1404 => x"0a",
  1405 => x"00",
  1406 => x"43",
  1407 => x"6f",
  1408 => x"6d",
  1409 => x"6d",
  1410 => x"61",
  1411 => x"6e",
  1412 => x"64",
  1413 => x"20",
  1414 => x"54",
  1415 => x"69",
  1416 => x"6d",
  1417 => x"65",
  1418 => x"6f",
  1419 => x"75",
  1420 => x"74",
  1421 => x"5f",
  1422 => x"45",
  1423 => x"72",
  1424 => x"72",
  1425 => x"6f",
  1426 => x"72",
  1427 => x"0d",
  1428 => x"0a",
  1429 => x"00",
  1430 => x"54",
  1431 => x"69",
  1432 => x"6d",
  1433 => x"65",
  1434 => x"6f",
  1435 => x"75",
  1436 => x"74",
  1437 => x"5f",
  1438 => x"45",
  1439 => x"72",
  1440 => x"72",
  1441 => x"6f",
  1442 => x"72",
  1443 => x"0d",
  1444 => x"0a",
  1445 => x"00",
  1446 => x"53",
  1447 => x"44",
  1448 => x"48",
  1449 => x"43",
  1450 => x"20",
  1451 => x"66",
  1452 => x"6f",
  1453 => x"75",
  1454 => x"6e",
  1455 => x"64",
  1456 => x"20",
  1457 => x"0d",
  1458 => x"0a",
  1459 => x"00",
  1460 => x"33",
  1461 => x"fc",
  1462 => x"ff",
  1463 => x"ff",
  1464 => x"00",
  1465 => x"7f",
  1466 => x"00",
  1467 => x"24",
  1468 => x"43",
  1469 => x"f9",
  1470 => x"81",
  1471 => x"00",
  1472 => x"00",
  1473 => x"00",
  1474 => x"33",
  1475 => x"7c",
  1476 => x"00",
  1477 => x"00",
  1478 => x"00",
  1479 => x"22",
  1480 => x"33",
  1481 => x"7c",
  1482 => x"00",
  1483 => x"96",
  1484 => x"00",
  1485 => x"1e",
  1486 => x"32",
  1487 => x"3c",
  1488 => x"00",
  1489 => x"c8",
  1490 => x"43",
  1491 => x"e9",
  1492 => x"00",
  1493 => x"20",
  1494 => x"33",
  1495 => x"7c",
  1496 => x"00",
  1497 => x"ff",
  1498 => x"00",
  1499 => x"24",
  1500 => x"51",
  1501 => x"c9",
  1502 => x"ff",
  1503 => x"f8",
  1504 => x"34",
  1505 => x"3c",
  1506 => x"00",
  1507 => x"32",
  1508 => x"61",
  1509 => x"00",
  1510 => x"fe",
  1511 => x"96",
  1512 => x"3f",
  1513 => x"69",
  1514 => x"00",
  1515 => x"24",
  1516 => x"ff",
  1517 => x"fe",
  1518 => x"33",
  1519 => x"7c",
  1520 => x"00",
  1521 => x"00",
  1522 => x"00",
  1523 => x"22",
  1524 => x"b0",
  1525 => x"3c",
  1526 => x"00",
  1527 => x"01",
  1528 => x"67",
  1529 => x"12",
  1530 => x"51",
  1531 => x"ca",
  1532 => x"ff",
  1533 => x"e8",
  1534 => x"48",
  1535 => x"7a",
  1536 => x"ff",
  1537 => x"6e",
  1538 => x"61",
  1539 => x"00",
  1540 => x"01",
  1541 => x"22",
  1542 => x"58",
  1543 => x"8f",
  1544 => x"70",
  1545 => x"ff",
  1546 => x"4e",
  1547 => x"75",
  1548 => x"22",
  1549 => x"3c",
  1550 => x"00",
  1551 => x"00",
  1552 => x"20",
  1553 => x"00",
  1554 => x"33",
  1555 => x"7c",
  1556 => x"00",
  1557 => x"ff",
  1558 => x"00",
  1559 => x"24",
  1560 => x"53",
  1561 => x"81",
  1562 => x"66",
  1563 => x"f6",
  1564 => x"61",
  1565 => x"00",
  1566 => x"fe",
  1567 => x"72",
  1568 => x"b0",
  1569 => x"3c",
  1570 => x"00",
  1571 => x"01",
  1572 => x"66",
  1573 => x"00",
  1574 => x"00",
  1575 => x"9e",
  1576 => x"33",
  1577 => x"7c",
  1578 => x"00",
  1579 => x"ff",
  1580 => x"00",
  1581 => x"24",
  1582 => x"33",
  1583 => x"7c",
  1584 => x"00",
  1585 => x"ff",
  1586 => x"00",
  1587 => x"24",
  1588 => x"33",
  1589 => x"7c",
  1590 => x"00",
  1591 => x"ff",
  1592 => x"00",
  1593 => x"24",
  1594 => x"30",
  1595 => x"29",
  1596 => x"00",
  1597 => x"24",
  1598 => x"0c",
  1599 => x"00",
  1600 => x"00",
  1601 => x"01",
  1602 => x"66",
  1603 => x"00",
  1604 => x"00",
  1605 => x"80",
  1606 => x"33",
  1607 => x"7c",
  1608 => x"00",
  1609 => x"ff",
  1610 => x"00",
  1611 => x"24",
  1612 => x"30",
  1613 => x"29",
  1614 => x"00",
  1615 => x"24",
  1616 => x"0c",
  1617 => x"00",
  1618 => x"00",
  1619 => x"aa",
  1620 => x"66",
  1621 => x"6e",
  1622 => x"3f",
  1623 => x"69",
  1624 => x"00",
  1625 => x"24",
  1626 => x"ff",
  1627 => x"fe",
  1628 => x"33",
  1629 => x"7c",
  1630 => x"00",
  1631 => x"00",
  1632 => x"00",
  1633 => x"22",
  1634 => x"48",
  1635 => x"7a",
  1636 => x"ff",
  1637 => x"42",
  1638 => x"61",
  1639 => x"00",
  1640 => x"00",
  1641 => x"be",
  1642 => x"58",
  1643 => x"8f",
  1644 => x"34",
  1645 => x"3c",
  1646 => x"00",
  1647 => x"32",
  1648 => x"53",
  1649 => x"42",
  1650 => x"67",
  1651 => x"50",
  1652 => x"32",
  1653 => x"3c",
  1654 => x"07",
  1655 => x"d0",
  1656 => x"33",
  1657 => x"7c",
  1658 => x"00",
  1659 => x"ff",
  1660 => x"00",
  1661 => x"24",
  1662 => x"51",
  1663 => x"c9",
  1664 => x"ff",
  1665 => x"f8",
  1666 => x"61",
  1667 => x"00",
  1668 => x"fe",
  1669 => x"28",
  1670 => x"b0",
  1671 => x"3c",
  1672 => x"00",
  1673 => x"01",
  1674 => x"66",
  1675 => x"e4",
  1676 => x"61",
  1677 => x"00",
  1678 => x"fe",
  1679 => x"10",
  1680 => x"66",
  1681 => x"de",
  1682 => x"61",
  1683 => x"00",
  1684 => x"fe",
  1685 => x"22",
  1686 => x"66",
  1687 => x"d8",
  1688 => x"33",
  1689 => x"7c",
  1690 => x"00",
  1691 => x"ff",
  1692 => x"00",
  1693 => x"24",
  1694 => x"30",
  1695 => x"29",
  1696 => x"00",
  1697 => x"24",
  1698 => x"c0",
  1699 => x"3c",
  1700 => x"00",
  1701 => x"40",
  1702 => x"66",
  1703 => x"08",
  1704 => x"33",
  1705 => x"fc",
  1706 => x"00",
  1707 => x"00",
  1708 => x"00",
  1709 => x"7f",
  1710 => x"00",
  1711 => x"24",
  1712 => x"33",
  1713 => x"7c",
  1714 => x"00",
  1715 => x"ff",
  1716 => x"00",
  1717 => x"24",
  1718 => x"33",
  1719 => x"7c",
  1720 => x"00",
  1721 => x"ff",
  1722 => x"00",
  1723 => x"24",
  1724 => x"33",
  1725 => x"7c",
  1726 => x"00",
  1727 => x"ff",
  1728 => x"00",
  1729 => x"24",
  1730 => x"60",
  1731 => x"3c",
  1732 => x"33",
  1733 => x"fc",
  1734 => x"00",
  1735 => x"00",
  1736 => x"00",
  1737 => x"7f",
  1738 => x"00",
  1739 => x"24",
  1740 => x"34",
  1741 => x"3c",
  1742 => x"00",
  1743 => x"0a",
  1744 => x"32",
  1745 => x"3c",
  1746 => x"07",
  1747 => x"d0",
  1748 => x"33",
  1749 => x"7c",
  1750 => x"00",
  1751 => x"ff",
  1752 => x"00",
  1753 => x"24",
  1754 => x"51",
  1755 => x"c9",
  1756 => x"ff",
  1757 => x"f8",
  1758 => x"61",
  1759 => x"00",
  1760 => x"fd",
  1761 => x"a6",
  1762 => x"67",
  1763 => x"1c",
  1764 => x"3f",
  1765 => x"69",
  1766 => x"00",
  1767 => x"24",
  1768 => x"ff",
  1769 => x"fe",
  1770 => x"33",
  1771 => x"7c",
  1772 => x"00",
  1773 => x"00",
  1774 => x"00",
  1775 => x"22",
  1776 => x"51",
  1777 => x"ca",
  1778 => x"ff",
  1779 => x"de",
  1780 => x"48",
  1781 => x"7a",
  1782 => x"fe",
  1783 => x"69",
  1784 => x"61",
  1785 => x"2c",
  1786 => x"58",
  1787 => x"8f",
  1788 => x"70",
  1789 => x"ff",
  1790 => x"4e",
  1791 => x"75",
  1792 => x"3f",
  1793 => x"69",
  1794 => x"00",
  1795 => x"24",
  1796 => x"ff",
  1797 => x"fe",
  1798 => x"33",
  1799 => x"7c",
  1800 => x"00",
  1801 => x"00",
  1802 => x"00",
  1803 => x"22",
  1804 => x"33",
  1805 => x"69",
  1806 => x"00",
  1807 => x"2c",
  1808 => x"00",
  1809 => x"1e",
  1810 => x"48",
  1811 => x"7a",
  1812 => x"fe",
  1813 => x"3f",
  1814 => x"61",
  1815 => x"0e",
  1816 => x"58",
  1817 => x"8f",
  1818 => x"33",
  1819 => x"fc",
  1820 => x"ff",
  1821 => x"ff",
  1822 => x"81",
  1823 => x"00",
  1824 => x"00",
  1825 => x"06",
  1826 => x"70",
  1827 => x"00",
  1828 => x"4e",
  1829 => x"75",
  1830 => x"2f",
  1831 => x"08",
  1832 => x"20",
  1833 => x"6f",
  1834 => x"00",
  1835 => x"08",
  1836 => x"61",
  1837 => x"04",
  1838 => x"20",
  1839 => x"5f",
  1840 => x"4e",
  1841 => x"75",
  1842 => x"48",
  1843 => x"e7",
  1844 => x"00",
  1845 => x"c0",
  1846 => x"22",
  1847 => x"39",
  1848 => x"00",
  1849 => x"7f",
  1850 => x"00",
  1851 => x"52",
  1852 => x"43",
  1853 => x"f9",
  1854 => x"80",
  1855 => x"00",
  1856 => x"08",
  1857 => x"00",
  1858 => x"10",
  1859 => x"18",
  1860 => x"67",
  1861 => x"08",
  1862 => x"13",
  1863 => x"80",
  1864 => x"10",
  1865 => x"00",
  1866 => x"52",
  1867 => x"41",
  1868 => x"60",
  1869 => x"f4",
  1870 => x"06",
  1871 => x"b9",
  1872 => x"00",
  1873 => x"00",
  1874 => x"00",
  1875 => x"4c",
  1876 => x"00",
  1877 => x"7f",
  1878 => x"00",
  1879 => x"52",
  1880 => x"4c",
  1881 => x"df",
  1882 => x"03",
  1883 => x"00",
  1884 => x"4e",
  1885 => x"75",
  1886 => x"4a",
  1887 => x"79",
  1888 => x"00",
  1889 => x"7f",
  1890 => x"00",
  1891 => x"24",
  1892 => x"67",
  1893 => x"1e",
  1894 => x"41",
  1895 => x"fa",
  1896 => x"00",
  1897 => x"08",
  1898 => x"48",
  1899 => x"7a",
  1900 => x"00",
  1901 => x"34",
  1902 => x"60",
  1903 => x"c2",
  1904 => x"53",
  1905 => x"44",
  1906 => x"48",
  1907 => x"43",
  1908 => x"20",
  1909 => x"66",
  1910 => x"6c",
  1911 => x"61",
  1912 => x"67",
  1913 => x"20",
  1914 => x"73",
  1915 => x"74",
  1916 => x"69",
  1917 => x"6c",
  1918 => x"6c",
  1919 => x"20",
  1920 => x"73",
  1921 => x"65",
  1922 => x"74",
  1923 => x"00",
  1924 => x"41",
  1925 => x"fa",
  1926 => x"00",
  1927 => x"08",
  1928 => x"48",
  1929 => x"7a",
  1930 => x"00",
  1931 => x"16",
  1932 => x"60",
  1933 => x"a4",
  1934 => x"53",
  1935 => x"44",
  1936 => x"48",
  1937 => x"43",
  1938 => x"20",
  1939 => x"66",
  1940 => x"6c",
  1941 => x"61",
  1942 => x"67",
  1943 => x"20",
  1944 => x"63",
  1945 => x"6c",
  1946 => x"65",
  1947 => x"61",
  1948 => x"72",
  1949 => x"65",
  1950 => x"64",
  1951 => x"00",
  1952 => x"61",
  1953 => x"00",
  1954 => x"02",
  1955 => x"0a",
  1956 => x"61",
  1957 => x"00",
  1958 => x"fc",
  1959 => x"46",
  1960 => x"66",
  1961 => x"46",
  1962 => x"2e",
  1963 => x"3c",
  1964 => x"00",
  1965 => x"00",
  1966 => x"01",
  1967 => x"ff",
  1968 => x"41",
  1969 => x"f9",
  1970 => x"00",
  1971 => x"7f",
  1972 => x"00",
  1973 => x"56",
  1974 => x"43",
  1975 => x"f9",
  1976 => x"80",
  1977 => x"00",
  1978 => x"08",
  1979 => x"00",
  1980 => x"10",
  1981 => x"18",
  1982 => x"12",
  1983 => x"c0",
  1984 => x"48",
  1985 => x"e7",
  1986 => x"01",
  1987 => x"c0",
  1988 => x"61",
  1989 => x"00",
  1990 => x"f9",
  1991 => x"70",
  1992 => x"4c",
  1993 => x"df",
  1994 => x"03",
  1995 => x"80",
  1996 => x"51",
  1997 => x"cf",
  1998 => x"ff",
  1999 => x"ee",
  2000 => x"20",
  2001 => x"39",
  2002 => x"00",
  2003 => x"7f",
  2004 => x"00",
  2005 => x"38",
  2006 => x"52",
  2007 => x"80",
  2008 => x"23",
  2009 => x"c0",
  2010 => x"00",
  2011 => x"7f",
  2012 => x"00",
  2013 => x"38",
  2014 => x"53",
  2015 => x"79",
  2016 => x"00",
  2017 => x"7f",
  2018 => x"00",
  2019 => x"36",
  2020 => x"66",
  2021 => x"be",
  2022 => x"61",
  2023 => x"00",
  2024 => x"02",
  2025 => x"7a",
  2026 => x"66",
  2027 => x"b4",
  2028 => x"20",
  2029 => x"08",
  2030 => x"4e",
  2031 => x"75",
  2032 => x"70",
  2033 => x"00",
  2034 => x"4e",
  2035 => x"75",
  2036 => x"33",
  2037 => x"fc",
  2038 => x"02",
  2039 => x"01",
  2040 => x"81",
  2041 => x"00",
  2042 => x"00",
  2043 => x"06",
  2044 => x"70",
  2045 => x"00",
  2046 => x"23",
  2047 => x"c0",
  2048 => x"00",
  2049 => x"7f",
  2050 => x"00",
  2051 => x"3e",
  2052 => x"33",
  2053 => x"fc",
  2054 => x"02",
  2055 => x"11",
  2056 => x"81",
  2057 => x"00",
  2058 => x"00",
  2059 => x"06",
  2060 => x"61",
  2061 => x"00",
  2062 => x"fb",
  2063 => x"de",
  2064 => x"66",
  2065 => x"5c",
  2066 => x"33",
  2067 => x"fc",
  2068 => x"02",
  2069 => x"02",
  2070 => x"81",
  2071 => x"00",
  2072 => x"00",
  2073 => x"06",
  2074 => x"0c",
  2075 => x"28",
  2076 => x"00",
  2077 => x"55",
  2078 => x"01",
  2079 => x"fe",
  2080 => x"66",
  2081 => x"4c",
  2082 => x"0c",
  2083 => x"28",
  2084 => x"00",
  2085 => x"aa",
  2086 => x"01",
  2087 => x"ff",
  2088 => x"66",
  2089 => x"44",
  2090 => x"30",
  2091 => x"39",
  2092 => x"00",
  2093 => x"7f",
  2094 => x"00",
  2095 => x"26",
  2096 => x"c0",
  2097 => x"7c",
  2098 => x"00",
  2099 => x"70",
  2100 => x"b0",
  2101 => x"7c",
  2102 => x"00",
  2103 => x"40",
  2104 => x"64",
  2105 => x"40",
  2106 => x"43",
  2107 => x"e8",
  2108 => x"01",
  2109 => x"be",
  2110 => x"d2",
  2111 => x"c0",
  2112 => x"33",
  2113 => x"fc",
  2114 => x"02",
  2115 => x"03",
  2116 => x"81",
  2117 => x"00",
  2118 => x"00",
  2119 => x"06",
  2120 => x"20",
  2121 => x"29",
  2122 => x"00",
  2123 => x"08",
  2124 => x"e0",
  2125 => x"58",
  2126 => x"48",
  2127 => x"40",
  2128 => x"e0",
  2129 => x"58",
  2130 => x"23",
  2131 => x"c0",
  2132 => x"00",
  2133 => x"7f",
  2134 => x"00",
  2135 => x"3e",
  2136 => x"61",
  2137 => x"00",
  2138 => x"fb",
  2139 => x"92",
  2140 => x"66",
  2141 => x"10",
  2142 => x"0c",
  2143 => x"28",
  2144 => x"00",
  2145 => x"55",
  2146 => x"01",
  2147 => x"fe",
  2148 => x"66",
  2149 => x"08",
  2150 => x"0c",
  2151 => x"28",
  2152 => x"00",
  2153 => x"aa",
  2154 => x"01",
  2155 => x"ff",
  2156 => x"67",
  2157 => x"0c",
  2158 => x"33",
  2159 => x"fc",
  2160 => x"f2",
  2161 => x"01",
  2162 => x"81",
  2163 => x"00",
  2164 => x"00",
  2165 => x"06",
  2166 => x"70",
  2167 => x"ff",
  2168 => x"4e",
  2169 => x"75",
  2170 => x"33",
  2171 => x"fc",
  2172 => x"02",
  2173 => x"04",
  2174 => x"81",
  2175 => x"00",
  2176 => x"00",
  2177 => x"06",
  2178 => x"0c",
  2179 => x"a8",
  2180 => x"46",
  2181 => x"41",
  2182 => x"54",
  2183 => x"31",
  2184 => x"00",
  2185 => x"36",
  2186 => x"66",
  2187 => x"24",
  2188 => x"13",
  2189 => x"fc",
  2190 => x"00",
  2191 => x"0c",
  2192 => x"00",
  2193 => x"7f",
  2194 => x"00",
  2195 => x"28",
  2196 => x"0c",
  2197 => x"a8",
  2198 => x"32",
  2199 => x"20",
  2200 => x"20",
  2201 => x"20",
  2202 => x"00",
  2203 => x"3a",
  2204 => x"67",
  2205 => x"36",
  2206 => x"13",
  2207 => x"fc",
  2208 => x"00",
  2209 => x"10",
  2210 => x"00",
  2211 => x"7f",
  2212 => x"00",
  2213 => x"28",
  2214 => x"0c",
  2215 => x"a8",
  2216 => x"36",
  2217 => x"20",
  2218 => x"20",
  2219 => x"20",
  2220 => x"00",
  2221 => x"3a",
  2222 => x"67",
  2223 => x"24",
  2224 => x"13",
  2225 => x"fc",
  2226 => x"00",
  2227 => x"00",
  2228 => x"00",
  2229 => x"7f",
  2230 => x"00",
  2231 => x"28",
  2232 => x"0c",
  2233 => x"a8",
  2234 => x"46",
  2235 => x"41",
  2236 => x"54",
  2237 => x"33",
  2238 => x"00",
  2239 => x"52",
  2240 => x"66",
  2241 => x"ac",
  2242 => x"0c",
  2243 => x"a8",
  2244 => x"32",
  2245 => x"20",
  2246 => x"20",
  2247 => x"20",
  2248 => x"00",
  2249 => x"56",
  2250 => x"66",
  2251 => x"a2",
  2252 => x"13",
  2253 => x"fc",
  2254 => x"00",
  2255 => x"20",
  2256 => x"00",
  2257 => x"7f",
  2258 => x"00",
  2259 => x"28",
  2260 => x"20",
  2261 => x"28",
  2262 => x"00",
  2263 => x"0a",
  2264 => x"c0",
  2265 => x"bc",
  2266 => x"00",
  2267 => x"ff",
  2268 => x"ff",
  2269 => x"00",
  2270 => x"0c",
  2271 => x"80",
  2272 => x"00",
  2273 => x"00",
  2274 => x"02",
  2275 => x"00",
  2276 => x"66",
  2277 => x"88",
  2278 => x"22",
  2279 => x"39",
  2280 => x"00",
  2281 => x"7f",
  2282 => x"00",
  2283 => x"3e",
  2284 => x"30",
  2285 => x"28",
  2286 => x"00",
  2287 => x"0e",
  2288 => x"e0",
  2289 => x"58",
  2290 => x"d2",
  2291 => x"80",
  2292 => x"23",
  2293 => x"c1",
  2294 => x"00",
  2295 => x"7f",
  2296 => x"00",
  2297 => x"42",
  2298 => x"0c",
  2299 => x"39",
  2300 => x"00",
  2301 => x"20",
  2302 => x"00",
  2303 => x"7f",
  2304 => x"00",
  2305 => x"28",
  2306 => x"66",
  2307 => x"24",
  2308 => x"20",
  2309 => x"28",
  2310 => x"00",
  2311 => x"2c",
  2312 => x"e0",
  2313 => x"58",
  2314 => x"48",
  2315 => x"40",
  2316 => x"e0",
  2317 => x"58",
  2318 => x"23",
  2319 => x"c0",
  2320 => x"00",
  2321 => x"7f",
  2322 => x"00",
  2323 => x"2a",
  2324 => x"20",
  2325 => x"28",
  2326 => x"00",
  2327 => x"24",
  2328 => x"e0",
  2329 => x"58",
  2330 => x"48",
  2331 => x"40",
  2332 => x"e0",
  2333 => x"58",
  2334 => x"d2",
  2335 => x"80",
  2336 => x"53",
  2337 => x"28",
  2338 => x"00",
  2339 => x"10",
  2340 => x"66",
  2341 => x"f8",
  2342 => x"60",
  2343 => x"32",
  2344 => x"70",
  2345 => x"00",
  2346 => x"23",
  2347 => x"c0",
  2348 => x"00",
  2349 => x"7f",
  2350 => x"00",
  2351 => x"2a",
  2352 => x"30",
  2353 => x"28",
  2354 => x"00",
  2355 => x"16",
  2356 => x"e0",
  2357 => x"58",
  2358 => x"d2",
  2359 => x"80",
  2360 => x"53",
  2361 => x"28",
  2362 => x"00",
  2363 => x"10",
  2364 => x"66",
  2365 => x"f8",
  2366 => x"23",
  2367 => x"c1",
  2368 => x"00",
  2369 => x"7f",
  2370 => x"00",
  2371 => x"2e",
  2372 => x"20",
  2373 => x"01",
  2374 => x"10",
  2375 => x"28",
  2376 => x"00",
  2377 => x"12",
  2378 => x"e1",
  2379 => x"48",
  2380 => x"10",
  2381 => x"28",
  2382 => x"00",
  2383 => x"11",
  2384 => x"33",
  2385 => x"c0",
  2386 => x"00",
  2387 => x"7f",
  2388 => x"00",
  2389 => x"4e",
  2390 => x"e8",
  2391 => x"48",
  2392 => x"d2",
  2393 => x"80",
  2394 => x"70",
  2395 => x"00",
  2396 => x"10",
  2397 => x"28",
  2398 => x"00",
  2399 => x"0d",
  2400 => x"33",
  2401 => x"c0",
  2402 => x"00",
  2403 => x"7f",
  2404 => x"00",
  2405 => x"4a",
  2406 => x"92",
  2407 => x"80",
  2408 => x"92",
  2409 => x"80",
  2410 => x"23",
  2411 => x"c1",
  2412 => x"00",
  2413 => x"7f",
  2414 => x"00",
  2415 => x"46",
  2416 => x"33",
  2417 => x"fc",
  2418 => x"02",
  2419 => x"05",
  2420 => x"81",
  2421 => x"00",
  2422 => x"00",
  2423 => x"06",
  2424 => x"70",
  2425 => x"00",
  2426 => x"4e",
  2427 => x"75",
  2428 => x"20",
  2429 => x"39",
  2430 => x"00",
  2431 => x"7f",
  2432 => x"00",
  2433 => x"2a",
  2434 => x"23",
  2435 => x"c0",
  2436 => x"00",
  2437 => x"7f",
  2438 => x"00",
  2439 => x"32",
  2440 => x"66",
  2441 => x"28",
  2442 => x"42",
  2443 => x"b9",
  2444 => x"00",
  2445 => x"7f",
  2446 => x"00",
  2447 => x"32",
  2448 => x"30",
  2449 => x"39",
  2450 => x"00",
  2451 => x"7f",
  2452 => x"00",
  2453 => x"4e",
  2454 => x"e8",
  2455 => x"48",
  2456 => x"33",
  2457 => x"c0",
  2458 => x"00",
  2459 => x"7f",
  2460 => x"00",
  2461 => x"36",
  2462 => x"20",
  2463 => x"39",
  2464 => x"00",
  2465 => x"7f",
  2466 => x"00",
  2467 => x"2e",
  2468 => x"23",
  2469 => x"c0",
  2470 => x"00",
  2471 => x"7f",
  2472 => x"00",
  2473 => x"38",
  2474 => x"4e",
  2475 => x"75",
  2476 => x"20",
  2477 => x"39",
  2478 => x"00",
  2479 => x"7f",
  2480 => x"00",
  2481 => x"32",
  2482 => x"32",
  2483 => x"39",
  2484 => x"00",
  2485 => x"7f",
  2486 => x"00",
  2487 => x"4a",
  2488 => x"33",
  2489 => x"c1",
  2490 => x"00",
  2491 => x"7f",
  2492 => x"00",
  2493 => x"36",
  2494 => x"e2",
  2495 => x"49",
  2496 => x"65",
  2497 => x"04",
  2498 => x"e3",
  2499 => x"88",
  2500 => x"60",
  2501 => x"f8",
  2502 => x"d0",
  2503 => x"b9",
  2504 => x"00",
  2505 => x"7f",
  2506 => x"00",
  2507 => x"46",
  2508 => x"23",
  2509 => x"c0",
  2510 => x"00",
  2511 => x"7f",
  2512 => x"00",
  2513 => x"38",
  2514 => x"4e",
  2515 => x"75",
  2516 => x"48",
  2517 => x"e7",
  2518 => x"20",
  2519 => x"20",
  2520 => x"24",
  2521 => x"49",
  2522 => x"61",
  2523 => x"00",
  2524 => x"fa",
  2525 => x"10",
  2526 => x"66",
  2527 => x"7a",
  2528 => x"74",
  2529 => x"0f",
  2530 => x"4a",
  2531 => x"10",
  2532 => x"67",
  2533 => x"74",
  2534 => x"70",
  2535 => x"0a",
  2536 => x"12",
  2537 => x"32",
  2538 => x"00",
  2539 => x"00",
  2540 => x"b2",
  2541 => x"30",
  2542 => x"00",
  2543 => x"00",
  2544 => x"67",
  2545 => x"0a",
  2546 => x"d2",
  2547 => x"3c",
  2548 => x"00",
  2549 => x"20",
  2550 => x"b2",
  2551 => x"30",
  2552 => x"00",
  2553 => x"00",
  2554 => x"66",
  2555 => x"36",
  2556 => x"51",
  2557 => x"c8",
  2558 => x"ff",
  2559 => x"ea",
  2560 => x"70",
  2561 => x"00",
  2562 => x"10",
  2563 => x"28",
  2564 => x"00",
  2565 => x"0b",
  2566 => x"33",
  2567 => x"c0",
  2568 => x"00",
  2569 => x"7f",
  2570 => x"00",
  2571 => x"3c",
  2572 => x"0c",
  2573 => x"39",
  2574 => x"00",
  2575 => x"20",
  2576 => x"00",
  2577 => x"7f",
  2578 => x"00",
  2579 => x"28",
  2580 => x"66",
  2581 => x"08",
  2582 => x"30",
  2583 => x"28",
  2584 => x"00",
  2585 => x"14",
  2586 => x"e0",
  2587 => x"58",
  2588 => x"48",
  2589 => x"40",
  2590 => x"30",
  2591 => x"28",
  2592 => x"00",
  2593 => x"1a",
  2594 => x"e0",
  2595 => x"58",
  2596 => x"23",
  2597 => x"c0",
  2598 => x"00",
  2599 => x"7f",
  2600 => x"00",
  2601 => x"32",
  2602 => x"4c",
  2603 => x"df",
  2604 => x"04",
  2605 => x"04",
  2606 => x"70",
  2607 => x"ff",
  2608 => x"4e",
  2609 => x"75",
  2610 => x"41",
  2611 => x"e8",
  2612 => x"00",
  2613 => x"20",
  2614 => x"51",
  2615 => x"ca",
  2616 => x"ff",
  2617 => x"aa",
  2618 => x"20",
  2619 => x"39",
  2620 => x"00",
  2621 => x"7f",
  2622 => x"00",
  2623 => x"38",
  2624 => x"52",
  2625 => x"80",
  2626 => x"23",
  2627 => x"c0",
  2628 => x"00",
  2629 => x"7f",
  2630 => x"00",
  2631 => x"38",
  2632 => x"53",
  2633 => x"79",
  2634 => x"00",
  2635 => x"7f",
  2636 => x"00",
  2637 => x"36",
  2638 => x"66",
  2639 => x"8a",
  2640 => x"61",
  2641 => x"10",
  2642 => x"67",
  2643 => x"06",
  2644 => x"61",
  2645 => x"00",
  2646 => x"ff",
  2647 => x"56",
  2648 => x"60",
  2649 => x"80",
  2650 => x"4c",
  2651 => x"df",
  2652 => x"04",
  2653 => x"04",
  2654 => x"70",
  2655 => x"00",
  2656 => x"4e",
  2657 => x"75",
  2658 => x"0c",
  2659 => x"39",
  2660 => x"00",
  2661 => x"20",
  2662 => x"00",
  2663 => x"7f",
  2664 => x"00",
  2665 => x"28",
  2666 => x"67",
  2667 => x"3e",
  2668 => x"0c",
  2669 => x"39",
  2670 => x"00",
  2671 => x"0c",
  2672 => x"00",
  2673 => x"7f",
  2674 => x"00",
  2675 => x"28",
  2676 => x"67",
  2677 => x"78",
  2678 => x"20",
  2679 => x"39",
  2680 => x"00",
  2681 => x"7f",
  2682 => x"00",
  2683 => x"32",
  2684 => x"e0",
  2685 => x"88",
  2686 => x"d0",
  2687 => x"b9",
  2688 => x"00",
  2689 => x"7f",
  2690 => x"00",
  2691 => x"42",
  2692 => x"61",
  2693 => x"00",
  2694 => x"f9",
  2695 => x"66",
  2696 => x"66",
  2697 => x"60",
  2698 => x"10",
  2699 => x"39",
  2700 => x"00",
  2701 => x"7f",
  2702 => x"00",
  2703 => x"35",
  2704 => x"d0",
  2705 => x"40",
  2706 => x"30",
  2707 => x"30",
  2708 => x"00",
  2709 => x"00",
  2710 => x"e0",
  2711 => x"58",
  2712 => x"23",
  2713 => x"c0",
  2714 => x"00",
  2715 => x"7f",
  2716 => x"00",
  2717 => x"32",
  2718 => x"80",
  2719 => x"bc",
  2720 => x"ff",
  2721 => x"ff",
  2722 => x"00",
  2723 => x"0f",
  2724 => x"b0",
  2725 => x"7c",
  2726 => x"ff",
  2727 => x"ff",
  2728 => x"4e",
  2729 => x"75",
  2730 => x"20",
  2731 => x"39",
  2732 => x"00",
  2733 => x"7f",
  2734 => x"00",
  2735 => x"32",
  2736 => x"ee",
  2737 => x"88",
  2738 => x"d0",
  2739 => x"b9",
  2740 => x"00",
  2741 => x"7f",
  2742 => x"00",
  2743 => x"42",
  2744 => x"61",
  2745 => x"00",
  2746 => x"f9",
  2747 => x"32",
  2748 => x"66",
  2749 => x"2c",
  2750 => x"10",
  2751 => x"39",
  2752 => x"00",
  2753 => x"7f",
  2754 => x"00",
  2755 => x"35",
  2756 => x"c0",
  2757 => x"7c",
  2758 => x"00",
  2759 => x"7f",
  2760 => x"d0",
  2761 => x"40",
  2762 => x"d0",
  2763 => x"40",
  2764 => x"20",
  2765 => x"30",
  2766 => x"00",
  2767 => x"00",
  2768 => x"e0",
  2769 => x"58",
  2770 => x"48",
  2771 => x"40",
  2772 => x"e0",
  2773 => x"58",
  2774 => x"23",
  2775 => x"c0",
  2776 => x"00",
  2777 => x"7f",
  2778 => x"00",
  2779 => x"32",
  2780 => x"80",
  2781 => x"bc",
  2782 => x"f0",
  2783 => x"00",
  2784 => x"00",
  2785 => x"07",
  2786 => x"b0",
  2787 => x"bc",
  2788 => x"ff",
  2789 => x"ff",
  2790 => x"ff",
  2791 => x"ff",
  2792 => x"4e",
  2793 => x"75",
  2794 => x"70",
  2795 => x"00",
  2796 => x"4e",
  2797 => x"75",
  2798 => x"2f",
  2799 => x"02",
  2800 => x"20",
  2801 => x"39",
  2802 => x"00",
  2803 => x"7f",
  2804 => x"00",
  2805 => x"32",
  2806 => x"22",
  2807 => x"00",
  2808 => x"d0",
  2809 => x"80",
  2810 => x"d0",
  2811 => x"81",
  2812 => x"22",
  2813 => x"00",
  2814 => x"e0",
  2815 => x"88",
  2816 => x"e4",
  2817 => x"88",
  2818 => x"d0",
  2819 => x"b9",
  2820 => x"00",
  2821 => x"7f",
  2822 => x"00",
  2823 => x"42",
  2824 => x"24",
  2825 => x"00",
  2826 => x"61",
  2827 => x"00",
  2828 => x"f8",
  2829 => x"e0",
  2830 => x"66",
  2831 => x"52",
  2832 => x"20",
  2833 => x"01",
  2834 => x"e2",
  2835 => x"88",
  2836 => x"c0",
  2837 => x"7c",
  2838 => x"01",
  2839 => x"ff",
  2840 => x"b0",
  2841 => x"7c",
  2842 => x"01",
  2843 => x"ff",
  2844 => x"66",
  2845 => x"14",
  2846 => x"10",
  2847 => x"30",
  2848 => x"00",
  2849 => x"00",
  2850 => x"c1",
  2851 => x"42",
  2852 => x"52",
  2853 => x"80",
  2854 => x"61",
  2855 => x"00",
  2856 => x"f8",
  2857 => x"c4",
  2858 => x"66",
  2859 => x"36",
  2860 => x"e1",
  2861 => x"4a",
  2862 => x"14",
  2863 => x"10",
  2864 => x"60",
  2865 => x"0a",
  2866 => x"14",
  2867 => x"30",
  2868 => x"00",
  2869 => x"00",
  2870 => x"e1",
  2871 => x"4a",
  2872 => x"14",
  2873 => x"30",
  2874 => x"00",
  2875 => x"01",
  2876 => x"e1",
  2877 => x"5a",
  2878 => x"c2",
  2879 => x"7c",
  2880 => x"00",
  2881 => x"01",
  2882 => x"67",
  2883 => x"02",
  2884 => x"e8",
  2885 => x"4a",
  2886 => x"c4",
  2887 => x"bc",
  2888 => x"00",
  2889 => x"00",
  2890 => x"0f",
  2891 => x"ff",
  2892 => x"23",
  2893 => x"c2",
  2894 => x"00",
  2895 => x"7f",
  2896 => x"00",
  2897 => x"32",
  2898 => x"84",
  2899 => x"bc",
  2900 => x"ff",
  2901 => x"ff",
  2902 => x"f0",
  2903 => x"0f",
  2904 => x"20",
  2905 => x"02",
  2906 => x"24",
  2907 => x"1f",
  2908 => x"b0",
  2909 => x"7c",
  2910 => x"ff",
  2911 => x"ff",
  2912 => x"4e",
  2913 => x"75",
  2914 => x"24",
  2915 => x"1f",
  2916 => x"70",
  2917 => x"00",
  2918 => x"4e",
  2919 => x"75",
  2920 => x"41",
  2921 => x"f9",
  2922 => x"00",
  2923 => x"7f",
  2924 => x"00",
  2925 => x"04",
  2926 => x"20",
  2927 => x"bc",
  2928 => x"12",
  2929 => x"34",
  2930 => x"56",
  2931 => x"78",
  2932 => x"21",
  2933 => x"7c",
  2934 => x"fe",
  2935 => x"dc",
  2936 => x"ba",
  2937 => x"98",
  2938 => x"00",
  2939 => x"04",
  2940 => x"21",
  2941 => x"7c",
  2942 => x"aa",
  2943 => x"55",
  2944 => x"cc",
  2945 => x"22",
  2946 => x"00",
  2947 => x"02",
  2948 => x"11",
  2949 => x"7c",
  2950 => x"00",
  2951 => x"33",
  2952 => x"00",
  2953 => x"03",
  2954 => x"11",
  2955 => x"7c",
  2956 => x"00",
  2957 => x"fe",
  2958 => x"00",
  2959 => x"04",
  2960 => x"20",
  2961 => x"10",
  2962 => x"22",
  2963 => x"28",
  2964 => x"00",
  2965 => x"04",
  2966 => x"90",
  2967 => x"bc",
  2968 => x"12",
  2969 => x"34",
  2970 => x"aa",
  2971 => x"33",
  2972 => x"92",
  2973 => x"bc",
  2974 => x"fe",
  2975 => x"22",
  2976 => x"ba",
  2977 => x"98",
  2978 => x"80",
  2979 => x"81",
  2980 => x"4e",
  2981 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


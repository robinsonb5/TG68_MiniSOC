library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"41",
    49 => x"fa",
    50 => x"00",
    51 => x"58",
    52 => x"61",
    53 => x"00",
    54 => x"02",
    55 => x"8c",
    56 => x"33",
    57 => x"fc",
    58 => x"0f",
    59 => x"00",
    60 => x"81",
    61 => x"00",
    62 => x"00",
    63 => x"06",
    64 => x"2e",
    65 => x"3c",
    66 => x"00",
    67 => x"00",
    68 => x"07",
    69 => x"ff",
    70 => x"41",
    71 => x"f9",
    72 => x"80",
    73 => x"00",
    74 => x"08",
    75 => x"00",
    76 => x"10",
    77 => x"fc",
    78 => x"00",
    79 => x"20",
    80 => x"51",
    81 => x"cf",
    82 => x"ff",
    83 => x"fa",
    84 => x"23",
    85 => x"fc",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"7f",
    92 => x"00",
    93 => x"52",
    94 => x"41",
    95 => x"fa",
    96 => x"00",
    97 => x"2a",
    98 => x"61",
    99 => x"00",
   100 => x"06",
   101 => x"6e",
   102 => x"61",
   103 => x"00",
   104 => x"02",
   105 => x"7a",
   106 => x"4b",
   107 => x"f9",
   108 => x"80",
   109 => x"00",
   110 => x"08",
   111 => x"00",
   112 => x"33",
   113 => x"fc",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"7f",
   118 => x"00",
   119 => x"0c",
   120 => x"30",
   121 => x"39",
   122 => x"81",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"08",
   127 => x"00",
   128 => x"00",
   129 => x"09",
   130 => x"67",
   131 => x"f4",
   132 => x"1a",
   133 => x"c0",
   134 => x"61",
   135 => x"4e",
   136 => x"60",
   137 => x"ee",
   138 => x"54",
   139 => x"65",
   140 => x"73",
   141 => x"74",
   142 => x"69",
   143 => x"6e",
   144 => x"67",
   145 => x"20",
   146 => x"73",
   147 => x"65",
   148 => x"72",
   149 => x"69",
   150 => x"61",
   151 => x"6c",
   152 => x"20",
   153 => x"6f",
   154 => x"75",
   155 => x"74",
   156 => x"70",
   157 => x"75",
   158 => x"74",
   159 => x"2e",
   160 => x"2e",
   161 => x"2e",
   162 => x"0d",
   163 => x"0a",
   164 => x"00",
   165 => x"00",
   166 => x"c0",
   167 => x"bc",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"df",
   172 => x"90",
   173 => x"3c",
   174 => x"00",
   175 => x"37",
   176 => x"6a",
   177 => x"04",
   178 => x"d0",
   179 => x"3c",
   180 => x"00",
   181 => x"27",
   182 => x"e9",
   183 => x"8e",
   184 => x"8c",
   185 => x"00",
   186 => x"20",
   187 => x"86",
   188 => x"4e",
   189 => x"75",
   190 => x"c0",
   191 => x"bc",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"df",
   196 => x"90",
   197 => x"3c",
   198 => x"00",
   199 => x"37",
   200 => x"6a",
   201 => x"04",
   202 => x"d0",
   203 => x"3c",
   204 => x"00",
   205 => x"27",
   206 => x"e9",
   207 => x"0f",
   208 => x"8e",
   209 => x"00",
   210 => x"10",
   211 => x"87",
   212 => x"4e",
   213 => x"75",
   214 => x"52",
   215 => x"79",
   216 => x"00",
   217 => x"7f",
   218 => x"00",
   219 => x"0c",
   220 => x"b0",
   221 => x"3c",
   222 => x"00",
   223 => x"53",
   224 => x"66",
   225 => x"2a",
   226 => x"33",
   227 => x"fc",
   228 => x"ff",
   229 => x"ff",
   230 => x"81",
   231 => x"00",
   232 => x"00",
   233 => x"06",
   234 => x"72",
   235 => x"00",
   236 => x"2e",
   237 => x"01",
   238 => x"2c",
   239 => x"01",
   240 => x"33",
   241 => x"c1",
   242 => x"00",
   243 => x"7f",
   244 => x"00",
   245 => x"0c",
   246 => x"23",
   247 => x"c1",
   248 => x"00",
   249 => x"7f",
   250 => x"00",
   251 => x"08",
   252 => x"23",
   253 => x"c1",
   254 => x"00",
   255 => x"7f",
   256 => x"00",
   257 => x"04",
   258 => x"23",
   259 => x"c1",
   260 => x"00",
   261 => x"7f",
   262 => x"00",
   263 => x"10",
   264 => x"60",
   265 => x"00",
   266 => x"01",
   267 => x"72",
   268 => x"2c",
   269 => x"39",
   270 => x"00",
   271 => x"7f",
   272 => x"00",
   273 => x"20",
   274 => x"2e",
   275 => x"39",
   276 => x"00",
   277 => x"7f",
   278 => x"00",
   279 => x"1c",
   280 => x"0c",
   281 => x"79",
   282 => x"00",
   283 => x"01",
   284 => x"00",
   285 => x"7f",
   286 => x"00",
   287 => x"0c",
   288 => x"66",
   289 => x"34",
   290 => x"33",
   291 => x"fc",
   292 => x"f0",
   293 => x"00",
   294 => x"81",
   295 => x"00",
   296 => x"00",
   297 => x"06",
   298 => x"41",
   299 => x"f9",
   300 => x"00",
   301 => x"7f",
   302 => x"00",
   303 => x"13",
   304 => x"61",
   305 => x"8c",
   306 => x"22",
   307 => x"39",
   308 => x"00",
   309 => x"7f",
   310 => x"00",
   311 => x"10",
   312 => x"b2",
   313 => x"bc",
   314 => x"00",
   315 => x"00",
   316 => x"00",
   317 => x"03",
   318 => x"6f",
   319 => x"08",
   320 => x"72",
   321 => x"0a",
   322 => x"92",
   323 => x"b9",
   324 => x"00",
   325 => x"7f",
   326 => x"00",
   327 => x"10",
   328 => x"52",
   329 => x"81",
   330 => x"e3",
   331 => x"89",
   332 => x"23",
   333 => x"c1",
   334 => x"00",
   335 => x"7f",
   336 => x"00",
   337 => x"14",
   338 => x"60",
   339 => x"00",
   340 => x"01",
   341 => x"28",
   342 => x"33",
   343 => x"f9",
   344 => x"00",
   345 => x"7f",
   346 => x"00",
   347 => x"12",
   348 => x"81",
   349 => x"00",
   350 => x"00",
   351 => x"06",
   352 => x"4a",
   353 => x"b9",
   354 => x"00",
   355 => x"7f",
   356 => x"00",
   357 => x"10",
   358 => x"67",
   359 => x"00",
   360 => x"01",
   361 => x"14",
   362 => x"0c",
   363 => x"b9",
   364 => x"00",
   365 => x"00",
   366 => x"00",
   367 => x"09",
   368 => x"00",
   369 => x"7f",
   370 => x"00",
   371 => x"10",
   372 => x"6e",
   373 => x"00",
   374 => x"00",
   375 => x"c0",
   376 => x"0c",
   377 => x"79",
   378 => x"00",
   379 => x"03",
   380 => x"00",
   381 => x"7f",
   382 => x"00",
   383 => x"0c",
   384 => x"6e",
   385 => x"16",
   386 => x"33",
   387 => x"fc",
   388 => x"0f",
   389 => x"00",
   390 => x"81",
   391 => x"00",
   392 => x"00",
   393 => x"06",
   394 => x"41",
   395 => x"f9",
   396 => x"00",
   397 => x"7f",
   398 => x"00",
   399 => x"07",
   400 => x"61",
   401 => x"00",
   402 => x"ff",
   403 => x"2c",
   404 => x"60",
   405 => x"00",
   406 => x"00",
   407 => x"e6",
   408 => x"22",
   409 => x"39",
   410 => x"00",
   411 => x"7f",
   412 => x"00",
   413 => x"14",
   414 => x"56",
   415 => x"41",
   416 => x"34",
   417 => x"39",
   418 => x"00",
   419 => x"7f",
   420 => x"00",
   421 => x"0c",
   422 => x"b4",
   423 => x"41",
   424 => x"6e",
   425 => x"20",
   426 => x"41",
   427 => x"f9",
   428 => x"00",
   429 => x"7f",
   430 => x"00",
   431 => x"08",
   432 => x"61",
   433 => x"00",
   434 => x"fe",
   435 => x"f4",
   436 => x"33",
   437 => x"f9",
   438 => x"00",
   439 => x"7f",
   440 => x"00",
   441 => x"0a",
   442 => x"81",
   443 => x"00",
   444 => x"00",
   445 => x"06",
   446 => x"33",
   447 => x"fc",
   448 => x"00",
   449 => x"01",
   450 => x"00",
   451 => x"7f",
   452 => x"00",
   453 => x"18",
   454 => x"60",
   455 => x"00",
   456 => x"00",
   457 => x"b4",
   458 => x"0c",
   459 => x"b9",
   460 => x"00",
   461 => x"00",
   462 => x"00",
   463 => x"03",
   464 => x"00",
   465 => x"7f",
   466 => x"00",
   467 => x"10",
   468 => x"6e",
   469 => x"60",
   470 => x"33",
   471 => x"fc",
   472 => x"00",
   473 => x"0f",
   474 => x"81",
   475 => x"00",
   476 => x"00",
   477 => x"06",
   478 => x"22",
   479 => x"39",
   480 => x"00",
   481 => x"7f",
   482 => x"00",
   483 => x"04",
   484 => x"e3",
   485 => x"89",
   486 => x"52",
   487 => x"81",
   488 => x"34",
   489 => x"39",
   490 => x"00",
   491 => x"7f",
   492 => x"00",
   493 => x"0c",
   494 => x"b4",
   495 => x"41",
   496 => x"6e",
   497 => x"2a",
   498 => x"20",
   499 => x"79",
   500 => x"00",
   501 => x"7f",
   502 => x"00",
   503 => x"08",
   504 => x"61",
   505 => x"00",
   506 => x"fe",
   507 => x"c4",
   508 => x"32",
   509 => x"39",
   510 => x"00",
   511 => x"7f",
   512 => x"00",
   513 => x"18",
   514 => x"53",
   515 => x"79",
   516 => x"00",
   517 => x"7f",
   518 => x"00",
   519 => x"18",
   520 => x"53",
   521 => x"41",
   522 => x"6a",
   523 => x"70",
   524 => x"52",
   525 => x"b9",
   526 => x"00",
   527 => x"7f",
   528 => x"00",
   529 => x"08",
   530 => x"33",
   531 => x"fc",
   532 => x"00",
   533 => x"01",
   534 => x"00",
   535 => x"7f",
   536 => x"00",
   537 => x"18",
   538 => x"60",
   539 => x"60",
   540 => x"30",
   541 => x"39",
   542 => x"00",
   543 => x"7f",
   544 => x"00",
   545 => x"18",
   546 => x"52",
   547 => x"40",
   548 => x"c0",
   549 => x"7c",
   550 => x"00",
   551 => x"01",
   552 => x"67",
   553 => x"52",
   554 => x"20",
   555 => x"79",
   556 => x"00",
   557 => x"7f",
   558 => x"00",
   559 => x"08",
   560 => x"e5",
   561 => x"88",
   562 => x"e1",
   563 => x"2f",
   564 => x"10",
   565 => x"87",
   566 => x"33",
   567 => x"fc",
   568 => x"f0",
   569 => x"f0",
   570 => x"81",
   571 => x"00",
   572 => x"00",
   573 => x"06",
   574 => x"0c",
   575 => x"b9",
   576 => x"00",
   577 => x"00",
   578 => x"00",
   579 => x"07",
   580 => x"00",
   581 => x"7f",
   582 => x"00",
   583 => x"10",
   584 => x"6d",
   585 => x"32",
   586 => x"33",
   587 => x"fc",
   588 => x"f0",
   589 => x"0f",
   590 => x"81",
   591 => x"00",
   592 => x"00",
   593 => x"06",
   594 => x"0c",
   595 => x"b9",
   596 => x"00",
   597 => x"00",
   598 => x"00",
   599 => x"09",
   600 => x"00",
   601 => x"7f",
   602 => x"00",
   603 => x"10",
   604 => x"6e",
   605 => x"1e",
   606 => x"33",
   607 => x"fc",
   608 => x"ff",
   609 => x"f0",
   610 => x"81",
   611 => x"00",
   612 => x"00",
   613 => x"06",
   614 => x"41",
   615 => x"fa",
   616 => x"00",
   617 => x"22",
   618 => x"61",
   619 => x"56",
   620 => x"2e",
   621 => x"b9",
   622 => x"00",
   623 => x"7f",
   624 => x"00",
   625 => x"08",
   626 => x"08",
   627 => x"b9",
   628 => x"00",
   629 => x"00",
   630 => x"81",
   631 => x"00",
   632 => x"00",
   633 => x"04",
   634 => x"4e",
   635 => x"75",
   636 => x"23",
   637 => x"c6",
   638 => x"00",
   639 => x"7f",
   640 => x"00",
   641 => x"20",
   642 => x"23",
   643 => x"c7",
   644 => x"00",
   645 => x"7f",
   646 => x"00",
   647 => x"1c",
   648 => x"4e",
   649 => x"75",
   650 => x"46",
   651 => x"69",
   652 => x"72",
   653 => x"6d",
   654 => x"77",
   655 => x"61",
   656 => x"72",
   657 => x"65",
   658 => x"20",
   659 => x"72",
   660 => x"65",
   661 => x"63",
   662 => x"65",
   663 => x"69",
   664 => x"76",
   665 => x"65",
   666 => x"64",
   667 => x"20",
   668 => x"2d",
   669 => x"20",
   670 => x"6c",
   671 => x"61",
   672 => x"75",
   673 => x"6e",
   674 => x"63",
   675 => x"68",
   676 => x"69",
   677 => x"6e",
   678 => x"67",
   679 => x"0d",
   680 => x"0a",
   681 => x"00",
   682 => x"48",
   683 => x"40",
   684 => x"30",
   685 => x"39",
   686 => x"81",
   687 => x"00",
   688 => x"00",
   689 => x"00",
   690 => x"08",
   691 => x"00",
   692 => x"00",
   693 => x"08",
   694 => x"67",
   695 => x"f4",
   696 => x"48",
   697 => x"40",
   698 => x"33",
   699 => x"c0",
   700 => x"81",
   701 => x"00",
   702 => x"00",
   703 => x"00",
   704 => x"4e",
   705 => x"75",
   706 => x"2f",
   707 => x"00",
   708 => x"70",
   709 => x"00",
   710 => x"30",
   711 => x"39",
   712 => x"81",
   713 => x"00",
   714 => x"00",
   715 => x"00",
   716 => x"08",
   717 => x"00",
   718 => x"00",
   719 => x"08",
   720 => x"67",
   721 => x"f4",
   722 => x"10",
   723 => x"18",
   724 => x"67",
   725 => x"08",
   726 => x"33",
   727 => x"c0",
   728 => x"81",
   729 => x"00",
   730 => x"00",
   731 => x"00",
   732 => x"60",
   733 => x"e8",
   734 => x"20",
   735 => x"1f",
   736 => x"4e",
   737 => x"75",
   738 => x"33",
   739 => x"fc",
   740 => x"00",
   741 => x"01",
   742 => x"81",
   743 => x"00",
   744 => x"00",
   745 => x"06",
   746 => x"41",
   747 => x"fa",
   748 => x"01",
   749 => x"fa",
   750 => x"61",
   751 => x"00",
   752 => x"03",
   753 => x"e2",
   754 => x"61",
   755 => x"00",
   756 => x"02",
   757 => x"60",
   758 => x"66",
   759 => x"5c",
   760 => x"33",
   761 => x"fc",
   762 => x"00",
   763 => x"02",
   764 => x"81",
   765 => x"00",
   766 => x"00",
   767 => x"06",
   768 => x"33",
   769 => x"fc",
   770 => x"00",
   771 => x"40",
   772 => x"00",
   773 => x"7f",
   774 => x"00",
   775 => x"26",
   776 => x"61",
   777 => x"00",
   778 => x"04",
   779 => x"8a",
   780 => x"67",
   781 => x"0c",
   782 => x"42",
   783 => x"79",
   784 => x"00",
   785 => x"7f",
   786 => x"00",
   787 => x"26",
   788 => x"61",
   789 => x"00",
   790 => x"04",
   791 => x"7e",
   792 => x"66",
   793 => x"28",
   794 => x"33",
   795 => x"fc",
   796 => x"00",
   797 => x"03",
   798 => x"81",
   799 => x"00",
   800 => x"00",
   801 => x"06",
   802 => x"61",
   803 => x"00",
   804 => x"05",
   805 => x"f8",
   806 => x"43",
   807 => x"fa",
   808 => x"00",
   809 => x"57",
   810 => x"61",
   811 => x"00",
   812 => x"06",
   813 => x"48",
   814 => x"67",
   815 => x"12",
   816 => x"41",
   817 => x"fa",
   818 => x"00",
   819 => x"47",
   820 => x"61",
   821 => x"00",
   822 => x"03",
   823 => x"9c",
   824 => x"30",
   825 => x"7c",
   826 => x"20",
   827 => x"00",
   828 => x"61",
   829 => x"00",
   830 => x"04",
   831 => x"02",
   832 => x"4e",
   833 => x"75",
   834 => x"33",
   835 => x"fc",
   836 => x"f0",
   837 => x"03",
   838 => x"81",
   839 => x"00",
   840 => x"00",
   841 => x"06",
   842 => x"41",
   843 => x"fa",
   844 => x"00",
   845 => x"29",
   846 => x"61",
   847 => x"00",
   848 => x"03",
   849 => x"82",
   850 => x"4e",
   851 => x"75",
   852 => x"33",
   853 => x"fc",
   854 => x"f0",
   855 => x"02",
   856 => x"81",
   857 => x"00",
   858 => x"00",
   859 => x"06",
   860 => x"41",
   861 => x"fa",
   862 => x"00",
   863 => x"08",
   864 => x"61",
   865 => x"00",
   866 => x"03",
   867 => x"70",
   868 => x"4e",
   869 => x"75",
   870 => x"53",
   871 => x"44",
   872 => x"20",
   873 => x"69",
   874 => x"6e",
   875 => x"69",
   876 => x"74",
   877 => x"20",
   878 => x"66",
   879 => x"61",
   880 => x"69",
   881 => x"6c",
   882 => x"65",
   883 => x"64",
   884 => x"00",
   885 => x"6e",
   886 => x"6f",
   887 => x"74",
   888 => x"20",
   889 => x"66",
   890 => x"6f",
   891 => x"75",
   892 => x"6e",
   893 => x"64",
   894 => x"20",
   895 => x"42",
   896 => x"4f",
   897 => x"4f",
   898 => x"54",
   899 => x"20",
   900 => x"20",
   901 => x"20",
   902 => x"20",
   903 => x"53",
   904 => x"52",
   905 => x"45",
   906 => x"00",
   907 => x"00",
   908 => x"33",
   909 => x"fc",
   910 => x"01",
   911 => x"00",
   912 => x"81",
   913 => x"00",
   914 => x"00",
   915 => x"06",
   916 => x"41",
   917 => x"f9",
   918 => x"00",
   919 => x"7f",
   920 => x"00",
   921 => x"56",
   922 => x"61",
   923 => x"00",
   924 => x"00",
   925 => x"c4",
   926 => x"66",
   927 => x"68",
   928 => x"33",
   929 => x"fc",
   930 => x"01",
   931 => x"01",
   932 => x"81",
   933 => x"00",
   934 => x"00",
   935 => x"06",
   936 => x"32",
   937 => x"3c",
   938 => x"4e",
   939 => x"20",
   940 => x"53",
   941 => x"41",
   942 => x"67",
   943 => x"44",
   944 => x"33",
   945 => x"fc",
   946 => x"01",
   947 => x"02",
   948 => x"81",
   949 => x"00",
   950 => x"00",
   951 => x"06",
   952 => x"33",
   953 => x"7c",
   954 => x"00",
   955 => x"ff",
   956 => x"00",
   957 => x"24",
   958 => x"30",
   959 => x"29",
   960 => x"00",
   961 => x"24",
   962 => x"b0",
   963 => x"3c",
   964 => x"00",
   965 => x"fe",
   966 => x"66",
   967 => x"e4",
   968 => x"30",
   969 => x"29",
   970 => x"01",
   971 => x"00",
   972 => x"32",
   973 => x"3c",
   974 => x"00",
   975 => x"7f",
   976 => x"20",
   977 => x"29",
   978 => x"01",
   979 => x"00",
   980 => x"20",
   981 => x"c0",
   982 => x"51",
   983 => x"c9",
   984 => x"ff",
   985 => x"f8",
   986 => x"30",
   987 => x"29",
   988 => x"00",
   989 => x"24",
   990 => x"33",
   991 => x"7c",
   992 => x"00",
   993 => x"00",
   994 => x"00",
   995 => x"22",
   996 => x"33",
   997 => x"fc",
   998 => x"01",
   999 => x"03",
  1000 => x"81",
  1001 => x"00",
  1002 => x"00",
  1003 => x"06",
  1004 => x"41",
  1005 => x"e8",
  1006 => x"fe",
  1007 => x"00",
  1008 => x"70",
  1009 => x"00",
  1010 => x"4e",
  1011 => x"75",
  1012 => x"33",
  1013 => x"fc",
  1014 => x"f1",
  1015 => x"02",
  1016 => x"81",
  1017 => x"00",
  1018 => x"00",
  1019 => x"06",
  1020 => x"41",
  1021 => x"fa",
  1022 => x"01",
  1023 => x"38",
  1024 => x"61",
  1025 => x"00",
  1026 => x"02",
  1027 => x"d0",
  1028 => x"70",
  1029 => x"fe",
  1030 => x"4e",
  1031 => x"75",
  1032 => x"33",
  1033 => x"fc",
  1034 => x"f1",
  1035 => x"03",
  1036 => x"81",
  1037 => x"00",
  1038 => x"00",
  1039 => x"06",
  1040 => x"41",
  1041 => x"fa",
  1042 => x"01",
  1043 => x"0c",
  1044 => x"61",
  1045 => x"00",
  1046 => x"02",
  1047 => x"bc",
  1048 => x"70",
  1049 => x"ff",
  1050 => x"4e",
  1051 => x"75",
  1052 => x"22",
  1053 => x"3c",
  1054 => x"00",
  1055 => x"95",
  1056 => x"00",
  1057 => x"40",
  1058 => x"70",
  1059 => x"00",
  1060 => x"60",
  1061 => x"40",
  1062 => x"22",
  1063 => x"3c",
  1064 => x"00",
  1065 => x"ff",
  1066 => x"00",
  1067 => x"41",
  1068 => x"70",
  1069 => x"00",
  1070 => x"60",
  1071 => x"36",
  1072 => x"22",
  1073 => x"3c",
  1074 => x"00",
  1075 => x"87",
  1076 => x"00",
  1077 => x"48",
  1078 => x"20",
  1079 => x"3c",
  1080 => x"00",
  1081 => x"00",
  1082 => x"01",
  1083 => x"aa",
  1084 => x"60",
  1085 => x"28",
  1086 => x"22",
  1087 => x"3c",
  1088 => x"00",
  1089 => x"87",
  1090 => x"00",
  1091 => x"69",
  1092 => x"20",
  1093 => x"3c",
  1094 => x"40",
  1095 => x"00",
  1096 => x"00",
  1097 => x"00",
  1098 => x"60",
  1099 => x"1a",
  1100 => x"22",
  1101 => x"3c",
  1102 => x"00",
  1103 => x"ff",
  1104 => x"00",
  1105 => x"77",
  1106 => x"70",
  1107 => x"00",
  1108 => x"60",
  1109 => x"10",
  1110 => x"22",
  1111 => x"3c",
  1112 => x"00",
  1113 => x"ff",
  1114 => x"00",
  1115 => x"7a",
  1116 => x"70",
  1117 => x"00",
  1118 => x"60",
  1119 => x"06",
  1120 => x"22",
  1121 => x"3c",
  1122 => x"00",
  1123 => x"ff",
  1124 => x"00",
  1125 => x"51",
  1126 => x"43",
  1127 => x"f9",
  1128 => x"81",
  1129 => x"00",
  1130 => x"00",
  1131 => x"00",
  1132 => x"33",
  1133 => x"7c",
  1134 => x"00",
  1135 => x"ff",
  1136 => x"00",
  1137 => x"24",
  1138 => x"3f",
  1139 => x"69",
  1140 => x"00",
  1141 => x"24",
  1142 => x"ff",
  1143 => x"fe",
  1144 => x"33",
  1145 => x"7c",
  1146 => x"00",
  1147 => x"01",
  1148 => x"00",
  1149 => x"22",
  1150 => x"33",
  1151 => x"7c",
  1152 => x"00",
  1153 => x"ff",
  1154 => x"00",
  1155 => x"24",
  1156 => x"33",
  1157 => x"41",
  1158 => x"00",
  1159 => x"24",
  1160 => x"48",
  1161 => x"41",
  1162 => x"4a",
  1163 => x"79",
  1164 => x"00",
  1165 => x"7f",
  1166 => x"00",
  1167 => x"24",
  1168 => x"67",
  1169 => x"16",
  1170 => x"e1",
  1171 => x"98",
  1172 => x"33",
  1173 => x"40",
  1174 => x"00",
  1175 => x"24",
  1176 => x"e1",
  1177 => x"98",
  1178 => x"33",
  1179 => x"40",
  1180 => x"00",
  1181 => x"24",
  1182 => x"e1",
  1183 => x"98",
  1184 => x"33",
  1185 => x"40",
  1186 => x"00",
  1187 => x"24",
  1188 => x"e1",
  1189 => x"98",
  1190 => x"60",
  1191 => x"18",
  1192 => x"d0",
  1193 => x"80",
  1194 => x"48",
  1195 => x"40",
  1196 => x"33",
  1197 => x"40",
  1198 => x"00",
  1199 => x"24",
  1200 => x"48",
  1201 => x"40",
  1202 => x"e1",
  1203 => x"58",
  1204 => x"33",
  1205 => x"40",
  1206 => x"00",
  1207 => x"24",
  1208 => x"e1",
  1209 => x"58",
  1210 => x"33",
  1211 => x"40",
  1212 => x"00",
  1213 => x"24",
  1214 => x"70",
  1215 => x"00",
  1216 => x"33",
  1217 => x"40",
  1218 => x"00",
  1219 => x"24",
  1220 => x"33",
  1221 => x"41",
  1222 => x"00",
  1223 => x"24",
  1224 => x"22",
  1225 => x"3c",
  1226 => x"00",
  1227 => x"00",
  1228 => x"01",
  1229 => x"90",
  1230 => x"53",
  1231 => x"81",
  1232 => x"67",
  1233 => x"10",
  1234 => x"33",
  1235 => x"7c",
  1236 => x"00",
  1237 => x"ff",
  1238 => x"00",
  1239 => x"24",
  1240 => x"30",
  1241 => x"29",
  1242 => x"00",
  1243 => x"24",
  1244 => x"b0",
  1245 => x"3c",
  1246 => x"00",
  1247 => x"ff",
  1248 => x"67",
  1249 => x"ec",
  1250 => x"80",
  1251 => x"00",
  1252 => x"4e",
  1253 => x"75",
  1254 => x"53",
  1255 => x"74",
  1256 => x"61",
  1257 => x"72",
  1258 => x"74",
  1259 => x"20",
  1260 => x"49",
  1261 => x"6e",
  1262 => x"69",
  1263 => x"74",
  1264 => x"0d",
  1265 => x"0a",
  1266 => x"00",
  1267 => x"49",
  1268 => x"6e",
  1269 => x"69",
  1270 => x"74",
  1271 => x"20",
  1272 => x"64",
  1273 => x"6f",
  1274 => x"6e",
  1275 => x"65",
  1276 => x"0d",
  1277 => x"0a",
  1278 => x"00",
  1279 => x"49",
  1280 => x"6e",
  1281 => x"69",
  1282 => x"74",
  1283 => x"20",
  1284 => x"66",
  1285 => x"61",
  1286 => x"69",
  1287 => x"6c",
  1288 => x"75",
  1289 => x"72",
  1290 => x"65",
  1291 => x"0d",
  1292 => x"0a",
  1293 => x"00",
  1294 => x"52",
  1295 => x"65",
  1296 => x"73",
  1297 => x"65",
  1298 => x"74",
  1299 => x"20",
  1300 => x"66",
  1301 => x"61",
  1302 => x"69",
  1303 => x"6c",
  1304 => x"75",
  1305 => x"72",
  1306 => x"65",
  1307 => x"0d",
  1308 => x"0a",
  1309 => x"00",
  1310 => x"43",
  1311 => x"6f",
  1312 => x"6d",
  1313 => x"6d",
  1314 => x"61",
  1315 => x"6e",
  1316 => x"64",
  1317 => x"20",
  1318 => x"54",
  1319 => x"69",
  1320 => x"6d",
  1321 => x"65",
  1322 => x"6f",
  1323 => x"75",
  1324 => x"74",
  1325 => x"5f",
  1326 => x"45",
  1327 => x"72",
  1328 => x"72",
  1329 => x"6f",
  1330 => x"72",
  1331 => x"0d",
  1332 => x"0a",
  1333 => x"00",
  1334 => x"54",
  1335 => x"69",
  1336 => x"6d",
  1337 => x"65",
  1338 => x"6f",
  1339 => x"75",
  1340 => x"74",
  1341 => x"5f",
  1342 => x"45",
  1343 => x"72",
  1344 => x"72",
  1345 => x"6f",
  1346 => x"72",
  1347 => x"0d",
  1348 => x"0a",
  1349 => x"00",
  1350 => x"53",
  1351 => x"44",
  1352 => x"48",
  1353 => x"43",
  1354 => x"20",
  1355 => x"66",
  1356 => x"6f",
  1357 => x"75",
  1358 => x"6e",
  1359 => x"64",
  1360 => x"20",
  1361 => x"0d",
  1362 => x"0a",
  1363 => x"00",
  1364 => x"33",
  1365 => x"fc",
  1366 => x"ff",
  1367 => x"ff",
  1368 => x"00",
  1369 => x"7f",
  1370 => x"00",
  1371 => x"24",
  1372 => x"43",
  1373 => x"f9",
  1374 => x"81",
  1375 => x"00",
  1376 => x"00",
  1377 => x"00",
  1378 => x"33",
  1379 => x"7c",
  1380 => x"00",
  1381 => x"00",
  1382 => x"00",
  1383 => x"22",
  1384 => x"33",
  1385 => x"7c",
  1386 => x"00",
  1387 => x"96",
  1388 => x"00",
  1389 => x"1e",
  1390 => x"32",
  1391 => x"3c",
  1392 => x"00",
  1393 => x"c8",
  1394 => x"43",
  1395 => x"e9",
  1396 => x"00",
  1397 => x"20",
  1398 => x"33",
  1399 => x"7c",
  1400 => x"00",
  1401 => x"ff",
  1402 => x"00",
  1403 => x"24",
  1404 => x"51",
  1405 => x"c9",
  1406 => x"ff",
  1407 => x"f8",
  1408 => x"34",
  1409 => x"3c",
  1410 => x"00",
  1411 => x"32",
  1412 => x"61",
  1413 => x"00",
  1414 => x"fe",
  1415 => x"96",
  1416 => x"3f",
  1417 => x"69",
  1418 => x"00",
  1419 => x"24",
  1420 => x"ff",
  1421 => x"fe",
  1422 => x"33",
  1423 => x"7c",
  1424 => x"00",
  1425 => x"00",
  1426 => x"00",
  1427 => x"22",
  1428 => x"b0",
  1429 => x"3c",
  1430 => x"00",
  1431 => x"01",
  1432 => x"67",
  1433 => x"12",
  1434 => x"51",
  1435 => x"ca",
  1436 => x"ff",
  1437 => x"e8",
  1438 => x"48",
  1439 => x"7a",
  1440 => x"ff",
  1441 => x"6e",
  1442 => x"61",
  1443 => x"00",
  1444 => x"01",
  1445 => x"22",
  1446 => x"58",
  1447 => x"8f",
  1448 => x"70",
  1449 => x"ff",
  1450 => x"4e",
  1451 => x"75",
  1452 => x"22",
  1453 => x"3c",
  1454 => x"00",
  1455 => x"00",
  1456 => x"20",
  1457 => x"00",
  1458 => x"33",
  1459 => x"7c",
  1460 => x"00",
  1461 => x"ff",
  1462 => x"00",
  1463 => x"24",
  1464 => x"53",
  1465 => x"81",
  1466 => x"66",
  1467 => x"f6",
  1468 => x"61",
  1469 => x"00",
  1470 => x"fe",
  1471 => x"72",
  1472 => x"b0",
  1473 => x"3c",
  1474 => x"00",
  1475 => x"01",
  1476 => x"66",
  1477 => x"00",
  1478 => x"00",
  1479 => x"9e",
  1480 => x"33",
  1481 => x"7c",
  1482 => x"00",
  1483 => x"ff",
  1484 => x"00",
  1485 => x"24",
  1486 => x"33",
  1487 => x"7c",
  1488 => x"00",
  1489 => x"ff",
  1490 => x"00",
  1491 => x"24",
  1492 => x"33",
  1493 => x"7c",
  1494 => x"00",
  1495 => x"ff",
  1496 => x"00",
  1497 => x"24",
  1498 => x"30",
  1499 => x"29",
  1500 => x"00",
  1501 => x"24",
  1502 => x"0c",
  1503 => x"00",
  1504 => x"00",
  1505 => x"01",
  1506 => x"66",
  1507 => x"00",
  1508 => x"00",
  1509 => x"80",
  1510 => x"33",
  1511 => x"7c",
  1512 => x"00",
  1513 => x"ff",
  1514 => x"00",
  1515 => x"24",
  1516 => x"30",
  1517 => x"29",
  1518 => x"00",
  1519 => x"24",
  1520 => x"0c",
  1521 => x"00",
  1522 => x"00",
  1523 => x"aa",
  1524 => x"66",
  1525 => x"6e",
  1526 => x"3f",
  1527 => x"69",
  1528 => x"00",
  1529 => x"24",
  1530 => x"ff",
  1531 => x"fe",
  1532 => x"33",
  1533 => x"7c",
  1534 => x"00",
  1535 => x"00",
  1536 => x"00",
  1537 => x"22",
  1538 => x"48",
  1539 => x"7a",
  1540 => x"ff",
  1541 => x"42",
  1542 => x"61",
  1543 => x"00",
  1544 => x"00",
  1545 => x"be",
  1546 => x"58",
  1547 => x"8f",
  1548 => x"34",
  1549 => x"3c",
  1550 => x"00",
  1551 => x"32",
  1552 => x"53",
  1553 => x"42",
  1554 => x"67",
  1555 => x"50",
  1556 => x"32",
  1557 => x"3c",
  1558 => x"07",
  1559 => x"d0",
  1560 => x"33",
  1561 => x"7c",
  1562 => x"00",
  1563 => x"ff",
  1564 => x"00",
  1565 => x"24",
  1566 => x"51",
  1567 => x"c9",
  1568 => x"ff",
  1569 => x"f8",
  1570 => x"61",
  1571 => x"00",
  1572 => x"fe",
  1573 => x"28",
  1574 => x"b0",
  1575 => x"3c",
  1576 => x"00",
  1577 => x"01",
  1578 => x"66",
  1579 => x"e4",
  1580 => x"61",
  1581 => x"00",
  1582 => x"fe",
  1583 => x"10",
  1584 => x"66",
  1585 => x"de",
  1586 => x"61",
  1587 => x"00",
  1588 => x"fe",
  1589 => x"22",
  1590 => x"66",
  1591 => x"d8",
  1592 => x"33",
  1593 => x"7c",
  1594 => x"00",
  1595 => x"ff",
  1596 => x"00",
  1597 => x"24",
  1598 => x"30",
  1599 => x"29",
  1600 => x"00",
  1601 => x"24",
  1602 => x"c0",
  1603 => x"3c",
  1604 => x"00",
  1605 => x"40",
  1606 => x"66",
  1607 => x"08",
  1608 => x"33",
  1609 => x"fc",
  1610 => x"00",
  1611 => x"00",
  1612 => x"00",
  1613 => x"7f",
  1614 => x"00",
  1615 => x"24",
  1616 => x"33",
  1617 => x"7c",
  1618 => x"00",
  1619 => x"ff",
  1620 => x"00",
  1621 => x"24",
  1622 => x"33",
  1623 => x"7c",
  1624 => x"00",
  1625 => x"ff",
  1626 => x"00",
  1627 => x"24",
  1628 => x"33",
  1629 => x"7c",
  1630 => x"00",
  1631 => x"ff",
  1632 => x"00",
  1633 => x"24",
  1634 => x"60",
  1635 => x"3c",
  1636 => x"33",
  1637 => x"fc",
  1638 => x"00",
  1639 => x"00",
  1640 => x"00",
  1641 => x"7f",
  1642 => x"00",
  1643 => x"24",
  1644 => x"34",
  1645 => x"3c",
  1646 => x"00",
  1647 => x"0a",
  1648 => x"32",
  1649 => x"3c",
  1650 => x"07",
  1651 => x"d0",
  1652 => x"33",
  1653 => x"7c",
  1654 => x"00",
  1655 => x"ff",
  1656 => x"00",
  1657 => x"24",
  1658 => x"51",
  1659 => x"c9",
  1660 => x"ff",
  1661 => x"f8",
  1662 => x"61",
  1663 => x"00",
  1664 => x"fd",
  1665 => x"a6",
  1666 => x"67",
  1667 => x"1c",
  1668 => x"3f",
  1669 => x"69",
  1670 => x"00",
  1671 => x"24",
  1672 => x"ff",
  1673 => x"fe",
  1674 => x"33",
  1675 => x"7c",
  1676 => x"00",
  1677 => x"00",
  1678 => x"00",
  1679 => x"22",
  1680 => x"51",
  1681 => x"ca",
  1682 => x"ff",
  1683 => x"de",
  1684 => x"48",
  1685 => x"7a",
  1686 => x"fe",
  1687 => x"69",
  1688 => x"61",
  1689 => x"2c",
  1690 => x"58",
  1691 => x"8f",
  1692 => x"70",
  1693 => x"ff",
  1694 => x"4e",
  1695 => x"75",
  1696 => x"3f",
  1697 => x"69",
  1698 => x"00",
  1699 => x"24",
  1700 => x"ff",
  1701 => x"fe",
  1702 => x"33",
  1703 => x"7c",
  1704 => x"00",
  1705 => x"00",
  1706 => x"00",
  1707 => x"22",
  1708 => x"33",
  1709 => x"69",
  1710 => x"00",
  1711 => x"2c",
  1712 => x"00",
  1713 => x"1e",
  1714 => x"48",
  1715 => x"7a",
  1716 => x"fe",
  1717 => x"3f",
  1718 => x"61",
  1719 => x"0e",
  1720 => x"58",
  1721 => x"8f",
  1722 => x"33",
  1723 => x"fc",
  1724 => x"ff",
  1725 => x"ff",
  1726 => x"81",
  1727 => x"00",
  1728 => x"00",
  1729 => x"06",
  1730 => x"70",
  1731 => x"00",
  1732 => x"4e",
  1733 => x"75",
  1734 => x"2f",
  1735 => x"08",
  1736 => x"20",
  1737 => x"6f",
  1738 => x"00",
  1739 => x"08",
  1740 => x"61",
  1741 => x"04",
  1742 => x"20",
  1743 => x"5f",
  1744 => x"4e",
  1745 => x"75",
  1746 => x"48",
  1747 => x"e7",
  1748 => x"00",
  1749 => x"c0",
  1750 => x"22",
  1751 => x"39",
  1752 => x"00",
  1753 => x"7f",
  1754 => x"00",
  1755 => x"52",
  1756 => x"43",
  1757 => x"f9",
  1758 => x"80",
  1759 => x"00",
  1760 => x"08",
  1761 => x"00",
  1762 => x"10",
  1763 => x"18",
  1764 => x"67",
  1765 => x"08",
  1766 => x"13",
  1767 => x"80",
  1768 => x"10",
  1769 => x"00",
  1770 => x"52",
  1771 => x"41",
  1772 => x"60",
  1773 => x"f4",
  1774 => x"06",
  1775 => x"b9",
  1776 => x"00",
  1777 => x"00",
  1778 => x"00",
  1779 => x"4c",
  1780 => x"00",
  1781 => x"7f",
  1782 => x"00",
  1783 => x"52",
  1784 => x"4c",
  1785 => x"df",
  1786 => x"03",
  1787 => x"00",
  1788 => x"4e",
  1789 => x"75",
  1790 => x"4a",
  1791 => x"79",
  1792 => x"00",
  1793 => x"7f",
  1794 => x"00",
  1795 => x"24",
  1796 => x"67",
  1797 => x"1e",
  1798 => x"41",
  1799 => x"fa",
  1800 => x"00",
  1801 => x"08",
  1802 => x"48",
  1803 => x"7a",
  1804 => x"00",
  1805 => x"34",
  1806 => x"60",
  1807 => x"c2",
  1808 => x"53",
  1809 => x"44",
  1810 => x"48",
  1811 => x"43",
  1812 => x"20",
  1813 => x"66",
  1814 => x"6c",
  1815 => x"61",
  1816 => x"67",
  1817 => x"20",
  1818 => x"73",
  1819 => x"74",
  1820 => x"69",
  1821 => x"6c",
  1822 => x"6c",
  1823 => x"20",
  1824 => x"73",
  1825 => x"65",
  1826 => x"74",
  1827 => x"00",
  1828 => x"41",
  1829 => x"fa",
  1830 => x"00",
  1831 => x"08",
  1832 => x"48",
  1833 => x"7a",
  1834 => x"00",
  1835 => x"16",
  1836 => x"60",
  1837 => x"a4",
  1838 => x"53",
  1839 => x"44",
  1840 => x"48",
  1841 => x"43",
  1842 => x"20",
  1843 => x"66",
  1844 => x"6c",
  1845 => x"61",
  1846 => x"67",
  1847 => x"20",
  1848 => x"63",
  1849 => x"6c",
  1850 => x"65",
  1851 => x"61",
  1852 => x"72",
  1853 => x"65",
  1854 => x"64",
  1855 => x"00",
  1856 => x"61",
  1857 => x"00",
  1858 => x"02",
  1859 => x"0a",
  1860 => x"61",
  1861 => x"00",
  1862 => x"fc",
  1863 => x"46",
  1864 => x"66",
  1865 => x"46",
  1866 => x"2e",
  1867 => x"3c",
  1868 => x"00",
  1869 => x"00",
  1870 => x"01",
  1871 => x"ff",
  1872 => x"41",
  1873 => x"f9",
  1874 => x"00",
  1875 => x"7f",
  1876 => x"00",
  1877 => x"56",
  1878 => x"43",
  1879 => x"f9",
  1880 => x"80",
  1881 => x"00",
  1882 => x"08",
  1883 => x"00",
  1884 => x"10",
  1885 => x"18",
  1886 => x"12",
  1887 => x"c0",
  1888 => x"48",
  1889 => x"e7",
  1890 => x"01",
  1891 => x"c0",
  1892 => x"61",
  1893 => x"00",
  1894 => x"f9",
  1895 => x"70",
  1896 => x"4c",
  1897 => x"df",
  1898 => x"03",
  1899 => x"80",
  1900 => x"51",
  1901 => x"cf",
  1902 => x"ff",
  1903 => x"ee",
  1904 => x"20",
  1905 => x"39",
  1906 => x"00",
  1907 => x"7f",
  1908 => x"00",
  1909 => x"38",
  1910 => x"52",
  1911 => x"80",
  1912 => x"23",
  1913 => x"c0",
  1914 => x"00",
  1915 => x"7f",
  1916 => x"00",
  1917 => x"38",
  1918 => x"53",
  1919 => x"79",
  1920 => x"00",
  1921 => x"7f",
  1922 => x"00",
  1923 => x"36",
  1924 => x"66",
  1925 => x"be",
  1926 => x"61",
  1927 => x"00",
  1928 => x"02",
  1929 => x"7a",
  1930 => x"66",
  1931 => x"b4",
  1932 => x"20",
  1933 => x"08",
  1934 => x"4e",
  1935 => x"75",
  1936 => x"70",
  1937 => x"00",
  1938 => x"4e",
  1939 => x"75",
  1940 => x"33",
  1941 => x"fc",
  1942 => x"02",
  1943 => x"01",
  1944 => x"81",
  1945 => x"00",
  1946 => x"00",
  1947 => x"06",
  1948 => x"70",
  1949 => x"00",
  1950 => x"23",
  1951 => x"c0",
  1952 => x"00",
  1953 => x"7f",
  1954 => x"00",
  1955 => x"3e",
  1956 => x"33",
  1957 => x"fc",
  1958 => x"02",
  1959 => x"11",
  1960 => x"81",
  1961 => x"00",
  1962 => x"00",
  1963 => x"06",
  1964 => x"61",
  1965 => x"00",
  1966 => x"fb",
  1967 => x"de",
  1968 => x"66",
  1969 => x"5c",
  1970 => x"33",
  1971 => x"fc",
  1972 => x"02",
  1973 => x"02",
  1974 => x"81",
  1975 => x"00",
  1976 => x"00",
  1977 => x"06",
  1978 => x"0c",
  1979 => x"28",
  1980 => x"00",
  1981 => x"55",
  1982 => x"01",
  1983 => x"fe",
  1984 => x"66",
  1985 => x"4c",
  1986 => x"0c",
  1987 => x"28",
  1988 => x"00",
  1989 => x"aa",
  1990 => x"01",
  1991 => x"ff",
  1992 => x"66",
  1993 => x"44",
  1994 => x"30",
  1995 => x"39",
  1996 => x"00",
  1997 => x"7f",
  1998 => x"00",
  1999 => x"26",
  2000 => x"c0",
  2001 => x"7c",
  2002 => x"00",
  2003 => x"70",
  2004 => x"b0",
  2005 => x"7c",
  2006 => x"00",
  2007 => x"40",
  2008 => x"64",
  2009 => x"40",
  2010 => x"43",
  2011 => x"e8",
  2012 => x"01",
  2013 => x"be",
  2014 => x"d2",
  2015 => x"c0",
  2016 => x"33",
  2017 => x"fc",
  2018 => x"02",
  2019 => x"03",
  2020 => x"81",
  2021 => x"00",
  2022 => x"00",
  2023 => x"06",
  2024 => x"20",
  2025 => x"29",
  2026 => x"00",
  2027 => x"08",
  2028 => x"e0",
  2029 => x"58",
  2030 => x"48",
  2031 => x"40",
  2032 => x"e0",
  2033 => x"58",
  2034 => x"23",
  2035 => x"c0",
  2036 => x"00",
  2037 => x"7f",
  2038 => x"00",
  2039 => x"3e",
  2040 => x"61",
  2041 => x"00",
  2042 => x"fb",
  2043 => x"92",
  2044 => x"66",
  2045 => x"10",
  2046 => x"0c",
  2047 => x"28",
  2048 => x"00",
  2049 => x"55",
  2050 => x"01",
  2051 => x"fe",
  2052 => x"66",
  2053 => x"08",
  2054 => x"0c",
  2055 => x"28",
  2056 => x"00",
  2057 => x"aa",
  2058 => x"01",
  2059 => x"ff",
  2060 => x"67",
  2061 => x"0c",
  2062 => x"33",
  2063 => x"fc",
  2064 => x"f2",
  2065 => x"01",
  2066 => x"81",
  2067 => x"00",
  2068 => x"00",
  2069 => x"06",
  2070 => x"70",
  2071 => x"ff",
  2072 => x"4e",
  2073 => x"75",
  2074 => x"33",
  2075 => x"fc",
  2076 => x"02",
  2077 => x"04",
  2078 => x"81",
  2079 => x"00",
  2080 => x"00",
  2081 => x"06",
  2082 => x"0c",
  2083 => x"a8",
  2084 => x"46",
  2085 => x"41",
  2086 => x"54",
  2087 => x"31",
  2088 => x"00",
  2089 => x"36",
  2090 => x"66",
  2091 => x"24",
  2092 => x"13",
  2093 => x"fc",
  2094 => x"00",
  2095 => x"0c",
  2096 => x"00",
  2097 => x"7f",
  2098 => x"00",
  2099 => x"28",
  2100 => x"0c",
  2101 => x"a8",
  2102 => x"32",
  2103 => x"20",
  2104 => x"20",
  2105 => x"20",
  2106 => x"00",
  2107 => x"3a",
  2108 => x"67",
  2109 => x"36",
  2110 => x"13",
  2111 => x"fc",
  2112 => x"00",
  2113 => x"10",
  2114 => x"00",
  2115 => x"7f",
  2116 => x"00",
  2117 => x"28",
  2118 => x"0c",
  2119 => x"a8",
  2120 => x"36",
  2121 => x"20",
  2122 => x"20",
  2123 => x"20",
  2124 => x"00",
  2125 => x"3a",
  2126 => x"67",
  2127 => x"24",
  2128 => x"13",
  2129 => x"fc",
  2130 => x"00",
  2131 => x"00",
  2132 => x"00",
  2133 => x"7f",
  2134 => x"00",
  2135 => x"28",
  2136 => x"0c",
  2137 => x"a8",
  2138 => x"46",
  2139 => x"41",
  2140 => x"54",
  2141 => x"33",
  2142 => x"00",
  2143 => x"52",
  2144 => x"66",
  2145 => x"ac",
  2146 => x"0c",
  2147 => x"a8",
  2148 => x"32",
  2149 => x"20",
  2150 => x"20",
  2151 => x"20",
  2152 => x"00",
  2153 => x"56",
  2154 => x"66",
  2155 => x"a2",
  2156 => x"13",
  2157 => x"fc",
  2158 => x"00",
  2159 => x"20",
  2160 => x"00",
  2161 => x"7f",
  2162 => x"00",
  2163 => x"28",
  2164 => x"20",
  2165 => x"28",
  2166 => x"00",
  2167 => x"0a",
  2168 => x"c0",
  2169 => x"bc",
  2170 => x"00",
  2171 => x"ff",
  2172 => x"ff",
  2173 => x"00",
  2174 => x"0c",
  2175 => x"80",
  2176 => x"00",
  2177 => x"00",
  2178 => x"02",
  2179 => x"00",
  2180 => x"66",
  2181 => x"88",
  2182 => x"22",
  2183 => x"39",
  2184 => x"00",
  2185 => x"7f",
  2186 => x"00",
  2187 => x"3e",
  2188 => x"30",
  2189 => x"28",
  2190 => x"00",
  2191 => x"0e",
  2192 => x"e0",
  2193 => x"58",
  2194 => x"d2",
  2195 => x"80",
  2196 => x"23",
  2197 => x"c1",
  2198 => x"00",
  2199 => x"7f",
  2200 => x"00",
  2201 => x"42",
  2202 => x"0c",
  2203 => x"39",
  2204 => x"00",
  2205 => x"20",
  2206 => x"00",
  2207 => x"7f",
  2208 => x"00",
  2209 => x"28",
  2210 => x"66",
  2211 => x"24",
  2212 => x"20",
  2213 => x"28",
  2214 => x"00",
  2215 => x"2c",
  2216 => x"e0",
  2217 => x"58",
  2218 => x"48",
  2219 => x"40",
  2220 => x"e0",
  2221 => x"58",
  2222 => x"23",
  2223 => x"c0",
  2224 => x"00",
  2225 => x"7f",
  2226 => x"00",
  2227 => x"2a",
  2228 => x"20",
  2229 => x"28",
  2230 => x"00",
  2231 => x"24",
  2232 => x"e0",
  2233 => x"58",
  2234 => x"48",
  2235 => x"40",
  2236 => x"e0",
  2237 => x"58",
  2238 => x"d2",
  2239 => x"80",
  2240 => x"53",
  2241 => x"28",
  2242 => x"00",
  2243 => x"10",
  2244 => x"66",
  2245 => x"f8",
  2246 => x"60",
  2247 => x"32",
  2248 => x"70",
  2249 => x"00",
  2250 => x"23",
  2251 => x"c0",
  2252 => x"00",
  2253 => x"7f",
  2254 => x"00",
  2255 => x"2a",
  2256 => x"30",
  2257 => x"28",
  2258 => x"00",
  2259 => x"16",
  2260 => x"e0",
  2261 => x"58",
  2262 => x"d2",
  2263 => x"80",
  2264 => x"53",
  2265 => x"28",
  2266 => x"00",
  2267 => x"10",
  2268 => x"66",
  2269 => x"f8",
  2270 => x"23",
  2271 => x"c1",
  2272 => x"00",
  2273 => x"7f",
  2274 => x"00",
  2275 => x"2e",
  2276 => x"20",
  2277 => x"01",
  2278 => x"10",
  2279 => x"28",
  2280 => x"00",
  2281 => x"12",
  2282 => x"e1",
  2283 => x"48",
  2284 => x"10",
  2285 => x"28",
  2286 => x"00",
  2287 => x"11",
  2288 => x"33",
  2289 => x"c0",
  2290 => x"00",
  2291 => x"7f",
  2292 => x"00",
  2293 => x"4e",
  2294 => x"e8",
  2295 => x"48",
  2296 => x"d2",
  2297 => x"80",
  2298 => x"70",
  2299 => x"00",
  2300 => x"10",
  2301 => x"28",
  2302 => x"00",
  2303 => x"0d",
  2304 => x"33",
  2305 => x"c0",
  2306 => x"00",
  2307 => x"7f",
  2308 => x"00",
  2309 => x"4a",
  2310 => x"92",
  2311 => x"80",
  2312 => x"92",
  2313 => x"80",
  2314 => x"23",
  2315 => x"c1",
  2316 => x"00",
  2317 => x"7f",
  2318 => x"00",
  2319 => x"46",
  2320 => x"33",
  2321 => x"fc",
  2322 => x"02",
  2323 => x"05",
  2324 => x"81",
  2325 => x"00",
  2326 => x"00",
  2327 => x"06",
  2328 => x"70",
  2329 => x"00",
  2330 => x"4e",
  2331 => x"75",
  2332 => x"20",
  2333 => x"39",
  2334 => x"00",
  2335 => x"7f",
  2336 => x"00",
  2337 => x"2a",
  2338 => x"23",
  2339 => x"c0",
  2340 => x"00",
  2341 => x"7f",
  2342 => x"00",
  2343 => x"32",
  2344 => x"66",
  2345 => x"28",
  2346 => x"42",
  2347 => x"b9",
  2348 => x"00",
  2349 => x"7f",
  2350 => x"00",
  2351 => x"32",
  2352 => x"30",
  2353 => x"39",
  2354 => x"00",
  2355 => x"7f",
  2356 => x"00",
  2357 => x"4e",
  2358 => x"e8",
  2359 => x"48",
  2360 => x"33",
  2361 => x"c0",
  2362 => x"00",
  2363 => x"7f",
  2364 => x"00",
  2365 => x"36",
  2366 => x"20",
  2367 => x"39",
  2368 => x"00",
  2369 => x"7f",
  2370 => x"00",
  2371 => x"2e",
  2372 => x"23",
  2373 => x"c0",
  2374 => x"00",
  2375 => x"7f",
  2376 => x"00",
  2377 => x"38",
  2378 => x"4e",
  2379 => x"75",
  2380 => x"20",
  2381 => x"39",
  2382 => x"00",
  2383 => x"7f",
  2384 => x"00",
  2385 => x"32",
  2386 => x"32",
  2387 => x"39",
  2388 => x"00",
  2389 => x"7f",
  2390 => x"00",
  2391 => x"4a",
  2392 => x"33",
  2393 => x"c1",
  2394 => x"00",
  2395 => x"7f",
  2396 => x"00",
  2397 => x"36",
  2398 => x"e2",
  2399 => x"49",
  2400 => x"65",
  2401 => x"04",
  2402 => x"e3",
  2403 => x"88",
  2404 => x"60",
  2405 => x"f8",
  2406 => x"d0",
  2407 => x"b9",
  2408 => x"00",
  2409 => x"7f",
  2410 => x"00",
  2411 => x"46",
  2412 => x"23",
  2413 => x"c0",
  2414 => x"00",
  2415 => x"7f",
  2416 => x"00",
  2417 => x"38",
  2418 => x"4e",
  2419 => x"75",
  2420 => x"48",
  2421 => x"e7",
  2422 => x"20",
  2423 => x"20",
  2424 => x"24",
  2425 => x"49",
  2426 => x"61",
  2427 => x"00",
  2428 => x"fa",
  2429 => x"10",
  2430 => x"66",
  2431 => x"7a",
  2432 => x"74",
  2433 => x"0f",
  2434 => x"4a",
  2435 => x"10",
  2436 => x"67",
  2437 => x"74",
  2438 => x"70",
  2439 => x"0a",
  2440 => x"12",
  2441 => x"32",
  2442 => x"00",
  2443 => x"00",
  2444 => x"b2",
  2445 => x"30",
  2446 => x"00",
  2447 => x"00",
  2448 => x"67",
  2449 => x"0a",
  2450 => x"d2",
  2451 => x"3c",
  2452 => x"00",
  2453 => x"20",
  2454 => x"b2",
  2455 => x"30",
  2456 => x"00",
  2457 => x"00",
  2458 => x"66",
  2459 => x"36",
  2460 => x"51",
  2461 => x"c8",
  2462 => x"ff",
  2463 => x"ea",
  2464 => x"70",
  2465 => x"00",
  2466 => x"10",
  2467 => x"28",
  2468 => x"00",
  2469 => x"0b",
  2470 => x"33",
  2471 => x"c0",
  2472 => x"00",
  2473 => x"7f",
  2474 => x"00",
  2475 => x"3c",
  2476 => x"0c",
  2477 => x"39",
  2478 => x"00",
  2479 => x"20",
  2480 => x"00",
  2481 => x"7f",
  2482 => x"00",
  2483 => x"28",
  2484 => x"66",
  2485 => x"08",
  2486 => x"30",
  2487 => x"28",
  2488 => x"00",
  2489 => x"14",
  2490 => x"e0",
  2491 => x"58",
  2492 => x"48",
  2493 => x"40",
  2494 => x"30",
  2495 => x"28",
  2496 => x"00",
  2497 => x"1a",
  2498 => x"e0",
  2499 => x"58",
  2500 => x"23",
  2501 => x"c0",
  2502 => x"00",
  2503 => x"7f",
  2504 => x"00",
  2505 => x"32",
  2506 => x"4c",
  2507 => x"df",
  2508 => x"04",
  2509 => x"04",
  2510 => x"70",
  2511 => x"ff",
  2512 => x"4e",
  2513 => x"75",
  2514 => x"41",
  2515 => x"e8",
  2516 => x"00",
  2517 => x"20",
  2518 => x"51",
  2519 => x"ca",
  2520 => x"ff",
  2521 => x"aa",
  2522 => x"20",
  2523 => x"39",
  2524 => x"00",
  2525 => x"7f",
  2526 => x"00",
  2527 => x"38",
  2528 => x"52",
  2529 => x"80",
  2530 => x"23",
  2531 => x"c0",
  2532 => x"00",
  2533 => x"7f",
  2534 => x"00",
  2535 => x"38",
  2536 => x"53",
  2537 => x"79",
  2538 => x"00",
  2539 => x"7f",
  2540 => x"00",
  2541 => x"36",
  2542 => x"66",
  2543 => x"8a",
  2544 => x"61",
  2545 => x"10",
  2546 => x"67",
  2547 => x"06",
  2548 => x"61",
  2549 => x"00",
  2550 => x"ff",
  2551 => x"56",
  2552 => x"60",
  2553 => x"80",
  2554 => x"4c",
  2555 => x"df",
  2556 => x"04",
  2557 => x"04",
  2558 => x"70",
  2559 => x"00",
  2560 => x"4e",
  2561 => x"75",
  2562 => x"0c",
  2563 => x"39",
  2564 => x"00",
  2565 => x"20",
  2566 => x"00",
  2567 => x"7f",
  2568 => x"00",
  2569 => x"28",
  2570 => x"67",
  2571 => x"3e",
  2572 => x"0c",
  2573 => x"39",
  2574 => x"00",
  2575 => x"0c",
  2576 => x"00",
  2577 => x"7f",
  2578 => x"00",
  2579 => x"28",
  2580 => x"67",
  2581 => x"78",
  2582 => x"20",
  2583 => x"39",
  2584 => x"00",
  2585 => x"7f",
  2586 => x"00",
  2587 => x"32",
  2588 => x"e0",
  2589 => x"88",
  2590 => x"d0",
  2591 => x"b9",
  2592 => x"00",
  2593 => x"7f",
  2594 => x"00",
  2595 => x"42",
  2596 => x"61",
  2597 => x"00",
  2598 => x"f9",
  2599 => x"66",
  2600 => x"66",
  2601 => x"60",
  2602 => x"10",
  2603 => x"39",
  2604 => x"00",
  2605 => x"7f",
  2606 => x"00",
  2607 => x"35",
  2608 => x"d0",
  2609 => x"40",
  2610 => x"30",
  2611 => x"30",
  2612 => x"00",
  2613 => x"00",
  2614 => x"e0",
  2615 => x"58",
  2616 => x"23",
  2617 => x"c0",
  2618 => x"00",
  2619 => x"7f",
  2620 => x"00",
  2621 => x"32",
  2622 => x"80",
  2623 => x"bc",
  2624 => x"ff",
  2625 => x"ff",
  2626 => x"00",
  2627 => x"0f",
  2628 => x"b0",
  2629 => x"7c",
  2630 => x"ff",
  2631 => x"ff",
  2632 => x"4e",
  2633 => x"75",
  2634 => x"20",
  2635 => x"39",
  2636 => x"00",
  2637 => x"7f",
  2638 => x"00",
  2639 => x"32",
  2640 => x"ee",
  2641 => x"88",
  2642 => x"d0",
  2643 => x"b9",
  2644 => x"00",
  2645 => x"7f",
  2646 => x"00",
  2647 => x"42",
  2648 => x"61",
  2649 => x"00",
  2650 => x"f9",
  2651 => x"32",
  2652 => x"66",
  2653 => x"2c",
  2654 => x"10",
  2655 => x"39",
  2656 => x"00",
  2657 => x"7f",
  2658 => x"00",
  2659 => x"35",
  2660 => x"c0",
  2661 => x"7c",
  2662 => x"00",
  2663 => x"7f",
  2664 => x"d0",
  2665 => x"40",
  2666 => x"d0",
  2667 => x"40",
  2668 => x"20",
  2669 => x"30",
  2670 => x"00",
  2671 => x"00",
  2672 => x"e0",
  2673 => x"58",
  2674 => x"48",
  2675 => x"40",
  2676 => x"e0",
  2677 => x"58",
  2678 => x"23",
  2679 => x"c0",
  2680 => x"00",
  2681 => x"7f",
  2682 => x"00",
  2683 => x"32",
  2684 => x"80",
  2685 => x"bc",
  2686 => x"f0",
  2687 => x"00",
  2688 => x"00",
  2689 => x"07",
  2690 => x"b0",
  2691 => x"bc",
  2692 => x"ff",
  2693 => x"ff",
  2694 => x"ff",
  2695 => x"ff",
  2696 => x"4e",
  2697 => x"75",
  2698 => x"70",
  2699 => x"00",
  2700 => x"4e",
  2701 => x"75",
  2702 => x"2f",
  2703 => x"02",
  2704 => x"20",
  2705 => x"39",
  2706 => x"00",
  2707 => x"7f",
  2708 => x"00",
  2709 => x"32",
  2710 => x"22",
  2711 => x"00",
  2712 => x"d0",
  2713 => x"80",
  2714 => x"d0",
  2715 => x"81",
  2716 => x"22",
  2717 => x"00",
  2718 => x"e0",
  2719 => x"88",
  2720 => x"e4",
  2721 => x"88",
  2722 => x"d0",
  2723 => x"b9",
  2724 => x"00",
  2725 => x"7f",
  2726 => x"00",
  2727 => x"42",
  2728 => x"24",
  2729 => x"00",
  2730 => x"61",
  2731 => x"00",
  2732 => x"f8",
  2733 => x"e0",
  2734 => x"66",
  2735 => x"52",
  2736 => x"20",
  2737 => x"01",
  2738 => x"e2",
  2739 => x"88",
  2740 => x"c0",
  2741 => x"7c",
  2742 => x"01",
  2743 => x"ff",
  2744 => x"b0",
  2745 => x"7c",
  2746 => x"01",
  2747 => x"ff",
  2748 => x"66",
  2749 => x"14",
  2750 => x"10",
  2751 => x"30",
  2752 => x"00",
  2753 => x"00",
  2754 => x"c1",
  2755 => x"42",
  2756 => x"52",
  2757 => x"80",
  2758 => x"61",
  2759 => x"00",
  2760 => x"f8",
  2761 => x"c4",
  2762 => x"66",
  2763 => x"36",
  2764 => x"e1",
  2765 => x"4a",
  2766 => x"14",
  2767 => x"10",
  2768 => x"60",
  2769 => x"0a",
  2770 => x"14",
  2771 => x"30",
  2772 => x"00",
  2773 => x"00",
  2774 => x"e1",
  2775 => x"4a",
  2776 => x"14",
  2777 => x"30",
  2778 => x"00",
  2779 => x"01",
  2780 => x"e1",
  2781 => x"5a",
  2782 => x"c2",
  2783 => x"7c",
  2784 => x"00",
  2785 => x"01",
  2786 => x"67",
  2787 => x"02",
  2788 => x"e8",
  2789 => x"4a",
  2790 => x"c4",
  2791 => x"bc",
  2792 => x"00",
  2793 => x"00",
  2794 => x"0f",
  2795 => x"ff",
  2796 => x"23",
  2797 => x"c2",
  2798 => x"00",
  2799 => x"7f",
  2800 => x"00",
  2801 => x"32",
  2802 => x"84",
  2803 => x"bc",
  2804 => x"ff",
  2805 => x"ff",
  2806 => x"f0",
  2807 => x"0f",
  2808 => x"20",
  2809 => x"02",
  2810 => x"24",
  2811 => x"1f",
  2812 => x"b0",
  2813 => x"7c",
  2814 => x"ff",
  2815 => x"ff",
  2816 => x"4e",
  2817 => x"75",
  2818 => x"24",
  2819 => x"1f",
  2820 => x"70",
  2821 => x"00",
  2822 => x"4e",
  2823 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


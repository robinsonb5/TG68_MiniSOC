library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"33",
    49 => x"fc",
    50 => x"00",
    51 => x"01",
    52 => x"81",
    53 => x"00",
    54 => x"00",
    55 => x"04",
    56 => x"41",
    57 => x"fa",
    58 => x"00",
    59 => x"74",
    60 => x"61",
    61 => x"00",
    62 => x"02",
    63 => x"d8",
    64 => x"33",
    65 => x"fc",
    66 => x"0f",
    67 => x"00",
    68 => x"81",
    69 => x"00",
    70 => x"00",
    71 => x"06",
    72 => x"2e",
    73 => x"3c",
    74 => x"00",
    75 => x"00",
    76 => x"07",
    77 => x"ff",
    78 => x"41",
    79 => x"f9",
    80 => x"80",
    81 => x"00",
    82 => x"08",
    83 => x"00",
    84 => x"10",
    85 => x"fc",
    86 => x"00",
    87 => x"20",
    88 => x"51",
    89 => x"cf",
    90 => x"ff",
    91 => x"fa",
    92 => x"23",
    93 => x"fc",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"7f",
   100 => x"00",
   101 => x"52",
   102 => x"41",
   103 => x"fa",
   104 => x"00",
   105 => x"46",
   106 => x"61",
   107 => x"00",
   108 => x"06",
   109 => x"ba",
   110 => x"61",
   111 => x"00",
   112 => x"0a",
   113 => x"ec",
   114 => x"4a",
   115 => x"80",
   116 => x"67",
   117 => x"0a",
   118 => x"41",
   119 => x"fa",
   120 => x"00",
   121 => x"6a",
   122 => x"61",
   123 => x"00",
   124 => x"06",
   125 => x"aa",
   126 => x"60",
   127 => x"fe",
   128 => x"41",
   129 => x"fa",
   130 => x"00",
   131 => x"49",
   132 => x"61",
   133 => x"00",
   134 => x"06",
   135 => x"a0",
   136 => x"61",
   137 => x"00",
   138 => x"02",
   139 => x"ac",
   140 => x"4b",
   141 => x"f9",
   142 => x"80",
   143 => x"00",
   144 => x"08",
   145 => x"00",
   146 => x"33",
   147 => x"fc",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"7f",
   152 => x"00",
   153 => x"0c",
   154 => x"30",
   155 => x"39",
   156 => x"81",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"08",
   161 => x"00",
   162 => x"00",
   163 => x"09",
   164 => x"67",
   165 => x"f4",
   166 => x"1a",
   167 => x"c0",
   168 => x"61",
   169 => x"00",
   170 => x"00",
   171 => x"80",
   172 => x"60",
   173 => x"ec",
   174 => x"43",
   175 => x"6f",
   176 => x"6e",
   177 => x"64",
   178 => x"75",
   179 => x"63",
   180 => x"74",
   181 => x"69",
   182 => x"6e",
   183 => x"67",
   184 => x"20",
   185 => x"73",
   186 => x"61",
   187 => x"6e",
   188 => x"69",
   189 => x"74",
   190 => x"79",
   191 => x"20",
   192 => x"63",
   193 => x"68",
   194 => x"65",
   195 => x"63",
   196 => x"6b",
   197 => x"2e",
   198 => x"2e",
   199 => x"2e",
   200 => x"0d",
   201 => x"0a",
   202 => x"00",
   203 => x"53",
   204 => x"61",
   205 => x"6e",
   206 => x"69",
   207 => x"74",
   208 => x"79",
   209 => x"20",
   210 => x"63",
   211 => x"68",
   212 => x"65",
   213 => x"63",
   214 => x"6b",
   215 => x"20",
   216 => x"70",
   217 => x"61",
   218 => x"73",
   219 => x"73",
   220 => x"65",
   221 => x"64",
   222 => x"2e",
   223 => x"0d",
   224 => x"0a",
   225 => x"00",
   226 => x"53",
   227 => x"61",
   228 => x"6e",
   229 => x"69",
   230 => x"74",
   231 => x"79",
   232 => x"20",
   233 => x"63",
   234 => x"68",
   235 => x"65",
   236 => x"63",
   237 => x"6b",
   238 => x"20",
   239 => x"66",
   240 => x"61",
   241 => x"69",
   242 => x"6c",
   243 => x"65",
   244 => x"64",
   245 => x"2e",
   246 => x"0d",
   247 => x"0a",
   248 => x"00",
   249 => x"00",
   250 => x"c0",
   251 => x"bc",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"df",
   256 => x"90",
   257 => x"3c",
   258 => x"00",
   259 => x"37",
   260 => x"6a",
   261 => x"04",
   262 => x"d0",
   263 => x"3c",
   264 => x"00",
   265 => x"27",
   266 => x"e9",
   267 => x"8e",
   268 => x"8c",
   269 => x"00",
   270 => x"20",
   271 => x"86",
   272 => x"4e",
   273 => x"75",
   274 => x"c0",
   275 => x"bc",
   276 => x"00",
   277 => x"00",
   278 => x"00",
   279 => x"df",
   280 => x"90",
   281 => x"3c",
   282 => x"00",
   283 => x"37",
   284 => x"6a",
   285 => x"04",
   286 => x"d0",
   287 => x"3c",
   288 => x"00",
   289 => x"27",
   290 => x"e9",
   291 => x"0f",
   292 => x"8e",
   293 => x"00",
   294 => x"10",
   295 => x"87",
   296 => x"4e",
   297 => x"75",
   298 => x"52",
   299 => x"79",
   300 => x"00",
   301 => x"7f",
   302 => x"00",
   303 => x"0c",
   304 => x"b0",
   305 => x"3c",
   306 => x"00",
   307 => x"53",
   308 => x"66",
   309 => x"2a",
   310 => x"33",
   311 => x"fc",
   312 => x"ff",
   313 => x"ff",
   314 => x"81",
   315 => x"00",
   316 => x"00",
   317 => x"06",
   318 => x"72",
   319 => x"00",
   320 => x"2e",
   321 => x"01",
   322 => x"2c",
   323 => x"01",
   324 => x"33",
   325 => x"c1",
   326 => x"00",
   327 => x"7f",
   328 => x"00",
   329 => x"0c",
   330 => x"23",
   331 => x"c1",
   332 => x"00",
   333 => x"7f",
   334 => x"00",
   335 => x"08",
   336 => x"23",
   337 => x"c1",
   338 => x"00",
   339 => x"7f",
   340 => x"00",
   341 => x"04",
   342 => x"23",
   343 => x"c1",
   344 => x"00",
   345 => x"7f",
   346 => x"00",
   347 => x"10",
   348 => x"60",
   349 => x"00",
   350 => x"01",
   351 => x"72",
   352 => x"2c",
   353 => x"39",
   354 => x"00",
   355 => x"7f",
   356 => x"00",
   357 => x"20",
   358 => x"2e",
   359 => x"39",
   360 => x"00",
   361 => x"7f",
   362 => x"00",
   363 => x"1c",
   364 => x"0c",
   365 => x"79",
   366 => x"00",
   367 => x"01",
   368 => x"00",
   369 => x"7f",
   370 => x"00",
   371 => x"0c",
   372 => x"66",
   373 => x"34",
   374 => x"33",
   375 => x"fc",
   376 => x"f0",
   377 => x"00",
   378 => x"81",
   379 => x"00",
   380 => x"00",
   381 => x"06",
   382 => x"41",
   383 => x"f9",
   384 => x"00",
   385 => x"7f",
   386 => x"00",
   387 => x"13",
   388 => x"61",
   389 => x"8c",
   390 => x"22",
   391 => x"39",
   392 => x"00",
   393 => x"7f",
   394 => x"00",
   395 => x"10",
   396 => x"b2",
   397 => x"bc",
   398 => x"00",
   399 => x"00",
   400 => x"00",
   401 => x"03",
   402 => x"6f",
   403 => x"08",
   404 => x"72",
   405 => x"0a",
   406 => x"92",
   407 => x"b9",
   408 => x"00",
   409 => x"7f",
   410 => x"00",
   411 => x"10",
   412 => x"52",
   413 => x"81",
   414 => x"e3",
   415 => x"89",
   416 => x"23",
   417 => x"c1",
   418 => x"00",
   419 => x"7f",
   420 => x"00",
   421 => x"14",
   422 => x"60",
   423 => x"00",
   424 => x"01",
   425 => x"28",
   426 => x"33",
   427 => x"f9",
   428 => x"00",
   429 => x"7f",
   430 => x"00",
   431 => x"12",
   432 => x"81",
   433 => x"00",
   434 => x"00",
   435 => x"06",
   436 => x"4a",
   437 => x"b9",
   438 => x"00",
   439 => x"7f",
   440 => x"00",
   441 => x"10",
   442 => x"67",
   443 => x"00",
   444 => x"01",
   445 => x"14",
   446 => x"0c",
   447 => x"b9",
   448 => x"00",
   449 => x"00",
   450 => x"00",
   451 => x"09",
   452 => x"00",
   453 => x"7f",
   454 => x"00",
   455 => x"10",
   456 => x"6e",
   457 => x"00",
   458 => x"00",
   459 => x"c0",
   460 => x"0c",
   461 => x"79",
   462 => x"00",
   463 => x"03",
   464 => x"00",
   465 => x"7f",
   466 => x"00",
   467 => x"0c",
   468 => x"6e",
   469 => x"16",
   470 => x"33",
   471 => x"fc",
   472 => x"0f",
   473 => x"00",
   474 => x"81",
   475 => x"00",
   476 => x"00",
   477 => x"06",
   478 => x"41",
   479 => x"f9",
   480 => x"00",
   481 => x"7f",
   482 => x"00",
   483 => x"07",
   484 => x"61",
   485 => x"00",
   486 => x"ff",
   487 => x"2c",
   488 => x"60",
   489 => x"00",
   490 => x"00",
   491 => x"e6",
   492 => x"22",
   493 => x"39",
   494 => x"00",
   495 => x"7f",
   496 => x"00",
   497 => x"14",
   498 => x"56",
   499 => x"41",
   500 => x"34",
   501 => x"39",
   502 => x"00",
   503 => x"7f",
   504 => x"00",
   505 => x"0c",
   506 => x"b4",
   507 => x"41",
   508 => x"6e",
   509 => x"20",
   510 => x"41",
   511 => x"f9",
   512 => x"00",
   513 => x"7f",
   514 => x"00",
   515 => x"08",
   516 => x"61",
   517 => x"00",
   518 => x"fe",
   519 => x"f4",
   520 => x"33",
   521 => x"f9",
   522 => x"00",
   523 => x"7f",
   524 => x"00",
   525 => x"0a",
   526 => x"81",
   527 => x"00",
   528 => x"00",
   529 => x"06",
   530 => x"33",
   531 => x"fc",
   532 => x"00",
   533 => x"01",
   534 => x"00",
   535 => x"7f",
   536 => x"00",
   537 => x"18",
   538 => x"60",
   539 => x"00",
   540 => x"00",
   541 => x"b4",
   542 => x"0c",
   543 => x"b9",
   544 => x"00",
   545 => x"00",
   546 => x"00",
   547 => x"03",
   548 => x"00",
   549 => x"7f",
   550 => x"00",
   551 => x"10",
   552 => x"6e",
   553 => x"60",
   554 => x"33",
   555 => x"fc",
   556 => x"00",
   557 => x"0f",
   558 => x"81",
   559 => x"00",
   560 => x"00",
   561 => x"06",
   562 => x"22",
   563 => x"39",
   564 => x"00",
   565 => x"7f",
   566 => x"00",
   567 => x"04",
   568 => x"e3",
   569 => x"89",
   570 => x"52",
   571 => x"81",
   572 => x"34",
   573 => x"39",
   574 => x"00",
   575 => x"7f",
   576 => x"00",
   577 => x"0c",
   578 => x"b4",
   579 => x"41",
   580 => x"6e",
   581 => x"2a",
   582 => x"20",
   583 => x"79",
   584 => x"00",
   585 => x"7f",
   586 => x"00",
   587 => x"08",
   588 => x"61",
   589 => x"00",
   590 => x"fe",
   591 => x"c4",
   592 => x"32",
   593 => x"39",
   594 => x"00",
   595 => x"7f",
   596 => x"00",
   597 => x"18",
   598 => x"53",
   599 => x"79",
   600 => x"00",
   601 => x"7f",
   602 => x"00",
   603 => x"18",
   604 => x"53",
   605 => x"41",
   606 => x"6a",
   607 => x"70",
   608 => x"52",
   609 => x"b9",
   610 => x"00",
   611 => x"7f",
   612 => x"00",
   613 => x"08",
   614 => x"33",
   615 => x"fc",
   616 => x"00",
   617 => x"01",
   618 => x"00",
   619 => x"7f",
   620 => x"00",
   621 => x"18",
   622 => x"60",
   623 => x"60",
   624 => x"30",
   625 => x"39",
   626 => x"00",
   627 => x"7f",
   628 => x"00",
   629 => x"18",
   630 => x"52",
   631 => x"40",
   632 => x"c0",
   633 => x"7c",
   634 => x"00",
   635 => x"01",
   636 => x"67",
   637 => x"52",
   638 => x"20",
   639 => x"79",
   640 => x"00",
   641 => x"7f",
   642 => x"00",
   643 => x"08",
   644 => x"e5",
   645 => x"88",
   646 => x"e1",
   647 => x"2f",
   648 => x"10",
   649 => x"87",
   650 => x"33",
   651 => x"fc",
   652 => x"f0",
   653 => x"f0",
   654 => x"81",
   655 => x"00",
   656 => x"00",
   657 => x"06",
   658 => x"0c",
   659 => x"b9",
   660 => x"00",
   661 => x"00",
   662 => x"00",
   663 => x"07",
   664 => x"00",
   665 => x"7f",
   666 => x"00",
   667 => x"10",
   668 => x"6d",
   669 => x"32",
   670 => x"33",
   671 => x"fc",
   672 => x"f0",
   673 => x"0f",
   674 => x"81",
   675 => x"00",
   676 => x"00",
   677 => x"06",
   678 => x"0c",
   679 => x"b9",
   680 => x"00",
   681 => x"00",
   682 => x"00",
   683 => x"09",
   684 => x"00",
   685 => x"7f",
   686 => x"00",
   687 => x"10",
   688 => x"6e",
   689 => x"1e",
   690 => x"33",
   691 => x"fc",
   692 => x"ff",
   693 => x"f0",
   694 => x"81",
   695 => x"00",
   696 => x"00",
   697 => x"06",
   698 => x"41",
   699 => x"fa",
   700 => x"00",
   701 => x"22",
   702 => x"61",
   703 => x"56",
   704 => x"2e",
   705 => x"b9",
   706 => x"00",
   707 => x"7f",
   708 => x"00",
   709 => x"08",
   710 => x"08",
   711 => x"b9",
   712 => x"00",
   713 => x"00",
   714 => x"81",
   715 => x"00",
   716 => x"00",
   717 => x"04",
   718 => x"4e",
   719 => x"75",
   720 => x"23",
   721 => x"c6",
   722 => x"00",
   723 => x"7f",
   724 => x"00",
   725 => x"20",
   726 => x"23",
   727 => x"c7",
   728 => x"00",
   729 => x"7f",
   730 => x"00",
   731 => x"1c",
   732 => x"4e",
   733 => x"75",
   734 => x"46",
   735 => x"69",
   736 => x"72",
   737 => x"6d",
   738 => x"77",
   739 => x"61",
   740 => x"72",
   741 => x"65",
   742 => x"20",
   743 => x"72",
   744 => x"65",
   745 => x"63",
   746 => x"65",
   747 => x"69",
   748 => x"76",
   749 => x"65",
   750 => x"64",
   751 => x"20",
   752 => x"2d",
   753 => x"20",
   754 => x"6c",
   755 => x"61",
   756 => x"75",
   757 => x"6e",
   758 => x"63",
   759 => x"68",
   760 => x"69",
   761 => x"6e",
   762 => x"67",
   763 => x"0d",
   764 => x"0a",
   765 => x"00",
   766 => x"48",
   767 => x"40",
   768 => x"30",
   769 => x"39",
   770 => x"81",
   771 => x"00",
   772 => x"00",
   773 => x"00",
   774 => x"08",
   775 => x"00",
   776 => x"00",
   777 => x"08",
   778 => x"67",
   779 => x"f4",
   780 => x"48",
   781 => x"40",
   782 => x"33",
   783 => x"c0",
   784 => x"81",
   785 => x"00",
   786 => x"00",
   787 => x"00",
   788 => x"4e",
   789 => x"75",
   790 => x"2f",
   791 => x"00",
   792 => x"70",
   793 => x"00",
   794 => x"30",
   795 => x"39",
   796 => x"81",
   797 => x"00",
   798 => x"00",
   799 => x"00",
   800 => x"08",
   801 => x"00",
   802 => x"00",
   803 => x"08",
   804 => x"67",
   805 => x"f4",
   806 => x"10",
   807 => x"18",
   808 => x"67",
   809 => x"08",
   810 => x"33",
   811 => x"c0",
   812 => x"81",
   813 => x"00",
   814 => x"00",
   815 => x"00",
   816 => x"60",
   817 => x"e8",
   818 => x"20",
   819 => x"1f",
   820 => x"4e",
   821 => x"75",
   822 => x"33",
   823 => x"fc",
   824 => x"00",
   825 => x"01",
   826 => x"81",
   827 => x"00",
   828 => x"00",
   829 => x"06",
   830 => x"41",
   831 => x"fa",
   832 => x"01",
   833 => x"fa",
   834 => x"61",
   835 => x"00",
   836 => x"03",
   837 => x"e2",
   838 => x"61",
   839 => x"00",
   840 => x"02",
   841 => x"60",
   842 => x"66",
   843 => x"5c",
   844 => x"33",
   845 => x"fc",
   846 => x"00",
   847 => x"02",
   848 => x"81",
   849 => x"00",
   850 => x"00",
   851 => x"06",
   852 => x"33",
   853 => x"fc",
   854 => x"00",
   855 => x"40",
   856 => x"00",
   857 => x"7f",
   858 => x"00",
   859 => x"26",
   860 => x"61",
   861 => x"00",
   862 => x"04",
   863 => x"8a",
   864 => x"67",
   865 => x"0c",
   866 => x"42",
   867 => x"79",
   868 => x"00",
   869 => x"7f",
   870 => x"00",
   871 => x"26",
   872 => x"61",
   873 => x"00",
   874 => x"04",
   875 => x"7e",
   876 => x"66",
   877 => x"28",
   878 => x"33",
   879 => x"fc",
   880 => x"00",
   881 => x"03",
   882 => x"81",
   883 => x"00",
   884 => x"00",
   885 => x"06",
   886 => x"61",
   887 => x"00",
   888 => x"05",
   889 => x"f8",
   890 => x"43",
   891 => x"fa",
   892 => x"00",
   893 => x"57",
   894 => x"61",
   895 => x"00",
   896 => x"06",
   897 => x"48",
   898 => x"67",
   899 => x"12",
   900 => x"41",
   901 => x"fa",
   902 => x"00",
   903 => x"47",
   904 => x"61",
   905 => x"00",
   906 => x"03",
   907 => x"9c",
   908 => x"30",
   909 => x"7c",
   910 => x"20",
   911 => x"00",
   912 => x"61",
   913 => x"00",
   914 => x"04",
   915 => x"02",
   916 => x"4e",
   917 => x"75",
   918 => x"33",
   919 => x"fc",
   920 => x"f0",
   921 => x"03",
   922 => x"81",
   923 => x"00",
   924 => x"00",
   925 => x"06",
   926 => x"41",
   927 => x"fa",
   928 => x"00",
   929 => x"29",
   930 => x"61",
   931 => x"00",
   932 => x"03",
   933 => x"82",
   934 => x"4e",
   935 => x"75",
   936 => x"33",
   937 => x"fc",
   938 => x"f0",
   939 => x"02",
   940 => x"81",
   941 => x"00",
   942 => x"00",
   943 => x"06",
   944 => x"41",
   945 => x"fa",
   946 => x"00",
   947 => x"08",
   948 => x"61",
   949 => x"00",
   950 => x"03",
   951 => x"70",
   952 => x"4e",
   953 => x"75",
   954 => x"53",
   955 => x"44",
   956 => x"20",
   957 => x"69",
   958 => x"6e",
   959 => x"69",
   960 => x"74",
   961 => x"20",
   962 => x"66",
   963 => x"61",
   964 => x"69",
   965 => x"6c",
   966 => x"65",
   967 => x"64",
   968 => x"00",
   969 => x"6e",
   970 => x"6f",
   971 => x"74",
   972 => x"20",
   973 => x"66",
   974 => x"6f",
   975 => x"75",
   976 => x"6e",
   977 => x"64",
   978 => x"20",
   979 => x"42",
   980 => x"4f",
   981 => x"4f",
   982 => x"54",
   983 => x"20",
   984 => x"20",
   985 => x"20",
   986 => x"20",
   987 => x"53",
   988 => x"52",
   989 => x"45",
   990 => x"00",
   991 => x"00",
   992 => x"33",
   993 => x"fc",
   994 => x"01",
   995 => x"00",
   996 => x"81",
   997 => x"00",
   998 => x"00",
   999 => x"06",
  1000 => x"41",
  1001 => x"f9",
  1002 => x"00",
  1003 => x"7f",
  1004 => x"00",
  1005 => x"56",
  1006 => x"61",
  1007 => x"00",
  1008 => x"00",
  1009 => x"c4",
  1010 => x"66",
  1011 => x"68",
  1012 => x"33",
  1013 => x"fc",
  1014 => x"01",
  1015 => x"01",
  1016 => x"81",
  1017 => x"00",
  1018 => x"00",
  1019 => x"06",
  1020 => x"32",
  1021 => x"3c",
  1022 => x"4e",
  1023 => x"20",
  1024 => x"53",
  1025 => x"41",
  1026 => x"67",
  1027 => x"44",
  1028 => x"33",
  1029 => x"fc",
  1030 => x"01",
  1031 => x"02",
  1032 => x"81",
  1033 => x"00",
  1034 => x"00",
  1035 => x"06",
  1036 => x"33",
  1037 => x"7c",
  1038 => x"00",
  1039 => x"ff",
  1040 => x"00",
  1041 => x"24",
  1042 => x"30",
  1043 => x"29",
  1044 => x"00",
  1045 => x"24",
  1046 => x"b0",
  1047 => x"3c",
  1048 => x"00",
  1049 => x"fe",
  1050 => x"66",
  1051 => x"e4",
  1052 => x"30",
  1053 => x"29",
  1054 => x"01",
  1055 => x"00",
  1056 => x"32",
  1057 => x"3c",
  1058 => x"00",
  1059 => x"7f",
  1060 => x"20",
  1061 => x"29",
  1062 => x"01",
  1063 => x"00",
  1064 => x"20",
  1065 => x"c0",
  1066 => x"51",
  1067 => x"c9",
  1068 => x"ff",
  1069 => x"f8",
  1070 => x"30",
  1071 => x"29",
  1072 => x"00",
  1073 => x"24",
  1074 => x"33",
  1075 => x"7c",
  1076 => x"00",
  1077 => x"00",
  1078 => x"00",
  1079 => x"22",
  1080 => x"33",
  1081 => x"fc",
  1082 => x"01",
  1083 => x"03",
  1084 => x"81",
  1085 => x"00",
  1086 => x"00",
  1087 => x"06",
  1088 => x"41",
  1089 => x"e8",
  1090 => x"fe",
  1091 => x"00",
  1092 => x"70",
  1093 => x"00",
  1094 => x"4e",
  1095 => x"75",
  1096 => x"33",
  1097 => x"fc",
  1098 => x"f1",
  1099 => x"02",
  1100 => x"81",
  1101 => x"00",
  1102 => x"00",
  1103 => x"06",
  1104 => x"41",
  1105 => x"fa",
  1106 => x"01",
  1107 => x"38",
  1108 => x"61",
  1109 => x"00",
  1110 => x"02",
  1111 => x"d0",
  1112 => x"70",
  1113 => x"fe",
  1114 => x"4e",
  1115 => x"75",
  1116 => x"33",
  1117 => x"fc",
  1118 => x"f1",
  1119 => x"03",
  1120 => x"81",
  1121 => x"00",
  1122 => x"00",
  1123 => x"06",
  1124 => x"41",
  1125 => x"fa",
  1126 => x"01",
  1127 => x"0c",
  1128 => x"61",
  1129 => x"00",
  1130 => x"02",
  1131 => x"bc",
  1132 => x"70",
  1133 => x"ff",
  1134 => x"4e",
  1135 => x"75",
  1136 => x"22",
  1137 => x"3c",
  1138 => x"00",
  1139 => x"95",
  1140 => x"00",
  1141 => x"40",
  1142 => x"70",
  1143 => x"00",
  1144 => x"60",
  1145 => x"40",
  1146 => x"22",
  1147 => x"3c",
  1148 => x"00",
  1149 => x"ff",
  1150 => x"00",
  1151 => x"41",
  1152 => x"70",
  1153 => x"00",
  1154 => x"60",
  1155 => x"36",
  1156 => x"22",
  1157 => x"3c",
  1158 => x"00",
  1159 => x"87",
  1160 => x"00",
  1161 => x"48",
  1162 => x"20",
  1163 => x"3c",
  1164 => x"00",
  1165 => x"00",
  1166 => x"01",
  1167 => x"aa",
  1168 => x"60",
  1169 => x"28",
  1170 => x"22",
  1171 => x"3c",
  1172 => x"00",
  1173 => x"87",
  1174 => x"00",
  1175 => x"69",
  1176 => x"20",
  1177 => x"3c",
  1178 => x"40",
  1179 => x"00",
  1180 => x"00",
  1181 => x"00",
  1182 => x"60",
  1183 => x"1a",
  1184 => x"22",
  1185 => x"3c",
  1186 => x"00",
  1187 => x"ff",
  1188 => x"00",
  1189 => x"77",
  1190 => x"70",
  1191 => x"00",
  1192 => x"60",
  1193 => x"10",
  1194 => x"22",
  1195 => x"3c",
  1196 => x"00",
  1197 => x"ff",
  1198 => x"00",
  1199 => x"7a",
  1200 => x"70",
  1201 => x"00",
  1202 => x"60",
  1203 => x"06",
  1204 => x"22",
  1205 => x"3c",
  1206 => x"00",
  1207 => x"ff",
  1208 => x"00",
  1209 => x"51",
  1210 => x"43",
  1211 => x"f9",
  1212 => x"81",
  1213 => x"00",
  1214 => x"00",
  1215 => x"00",
  1216 => x"33",
  1217 => x"7c",
  1218 => x"00",
  1219 => x"ff",
  1220 => x"00",
  1221 => x"24",
  1222 => x"3f",
  1223 => x"69",
  1224 => x"00",
  1225 => x"24",
  1226 => x"ff",
  1227 => x"fe",
  1228 => x"33",
  1229 => x"7c",
  1230 => x"00",
  1231 => x"01",
  1232 => x"00",
  1233 => x"22",
  1234 => x"33",
  1235 => x"7c",
  1236 => x"00",
  1237 => x"ff",
  1238 => x"00",
  1239 => x"24",
  1240 => x"33",
  1241 => x"41",
  1242 => x"00",
  1243 => x"24",
  1244 => x"48",
  1245 => x"41",
  1246 => x"4a",
  1247 => x"79",
  1248 => x"00",
  1249 => x"7f",
  1250 => x"00",
  1251 => x"24",
  1252 => x"67",
  1253 => x"16",
  1254 => x"e1",
  1255 => x"98",
  1256 => x"33",
  1257 => x"40",
  1258 => x"00",
  1259 => x"24",
  1260 => x"e1",
  1261 => x"98",
  1262 => x"33",
  1263 => x"40",
  1264 => x"00",
  1265 => x"24",
  1266 => x"e1",
  1267 => x"98",
  1268 => x"33",
  1269 => x"40",
  1270 => x"00",
  1271 => x"24",
  1272 => x"e1",
  1273 => x"98",
  1274 => x"60",
  1275 => x"18",
  1276 => x"d0",
  1277 => x"80",
  1278 => x"48",
  1279 => x"40",
  1280 => x"33",
  1281 => x"40",
  1282 => x"00",
  1283 => x"24",
  1284 => x"48",
  1285 => x"40",
  1286 => x"e1",
  1287 => x"58",
  1288 => x"33",
  1289 => x"40",
  1290 => x"00",
  1291 => x"24",
  1292 => x"e1",
  1293 => x"58",
  1294 => x"33",
  1295 => x"40",
  1296 => x"00",
  1297 => x"24",
  1298 => x"70",
  1299 => x"00",
  1300 => x"33",
  1301 => x"40",
  1302 => x"00",
  1303 => x"24",
  1304 => x"33",
  1305 => x"41",
  1306 => x"00",
  1307 => x"24",
  1308 => x"22",
  1309 => x"3c",
  1310 => x"00",
  1311 => x"00",
  1312 => x"01",
  1313 => x"90",
  1314 => x"53",
  1315 => x"81",
  1316 => x"67",
  1317 => x"10",
  1318 => x"33",
  1319 => x"7c",
  1320 => x"00",
  1321 => x"ff",
  1322 => x"00",
  1323 => x"24",
  1324 => x"30",
  1325 => x"29",
  1326 => x"00",
  1327 => x"24",
  1328 => x"b0",
  1329 => x"3c",
  1330 => x"00",
  1331 => x"ff",
  1332 => x"67",
  1333 => x"ec",
  1334 => x"80",
  1335 => x"00",
  1336 => x"4e",
  1337 => x"75",
  1338 => x"53",
  1339 => x"74",
  1340 => x"61",
  1341 => x"72",
  1342 => x"74",
  1343 => x"20",
  1344 => x"49",
  1345 => x"6e",
  1346 => x"69",
  1347 => x"74",
  1348 => x"0d",
  1349 => x"0a",
  1350 => x"00",
  1351 => x"49",
  1352 => x"6e",
  1353 => x"69",
  1354 => x"74",
  1355 => x"20",
  1356 => x"64",
  1357 => x"6f",
  1358 => x"6e",
  1359 => x"65",
  1360 => x"0d",
  1361 => x"0a",
  1362 => x"00",
  1363 => x"49",
  1364 => x"6e",
  1365 => x"69",
  1366 => x"74",
  1367 => x"20",
  1368 => x"66",
  1369 => x"61",
  1370 => x"69",
  1371 => x"6c",
  1372 => x"75",
  1373 => x"72",
  1374 => x"65",
  1375 => x"0d",
  1376 => x"0a",
  1377 => x"00",
  1378 => x"52",
  1379 => x"65",
  1380 => x"73",
  1381 => x"65",
  1382 => x"74",
  1383 => x"20",
  1384 => x"66",
  1385 => x"61",
  1386 => x"69",
  1387 => x"6c",
  1388 => x"75",
  1389 => x"72",
  1390 => x"65",
  1391 => x"0d",
  1392 => x"0a",
  1393 => x"00",
  1394 => x"43",
  1395 => x"6f",
  1396 => x"6d",
  1397 => x"6d",
  1398 => x"61",
  1399 => x"6e",
  1400 => x"64",
  1401 => x"20",
  1402 => x"54",
  1403 => x"69",
  1404 => x"6d",
  1405 => x"65",
  1406 => x"6f",
  1407 => x"75",
  1408 => x"74",
  1409 => x"5f",
  1410 => x"45",
  1411 => x"72",
  1412 => x"72",
  1413 => x"6f",
  1414 => x"72",
  1415 => x"0d",
  1416 => x"0a",
  1417 => x"00",
  1418 => x"54",
  1419 => x"69",
  1420 => x"6d",
  1421 => x"65",
  1422 => x"6f",
  1423 => x"75",
  1424 => x"74",
  1425 => x"5f",
  1426 => x"45",
  1427 => x"72",
  1428 => x"72",
  1429 => x"6f",
  1430 => x"72",
  1431 => x"0d",
  1432 => x"0a",
  1433 => x"00",
  1434 => x"53",
  1435 => x"44",
  1436 => x"48",
  1437 => x"43",
  1438 => x"20",
  1439 => x"66",
  1440 => x"6f",
  1441 => x"75",
  1442 => x"6e",
  1443 => x"64",
  1444 => x"20",
  1445 => x"0d",
  1446 => x"0a",
  1447 => x"00",
  1448 => x"33",
  1449 => x"fc",
  1450 => x"ff",
  1451 => x"ff",
  1452 => x"00",
  1453 => x"7f",
  1454 => x"00",
  1455 => x"24",
  1456 => x"43",
  1457 => x"f9",
  1458 => x"81",
  1459 => x"00",
  1460 => x"00",
  1461 => x"00",
  1462 => x"33",
  1463 => x"7c",
  1464 => x"00",
  1465 => x"00",
  1466 => x"00",
  1467 => x"22",
  1468 => x"33",
  1469 => x"7c",
  1470 => x"00",
  1471 => x"96",
  1472 => x"00",
  1473 => x"1e",
  1474 => x"32",
  1475 => x"3c",
  1476 => x"00",
  1477 => x"c8",
  1478 => x"43",
  1479 => x"e9",
  1480 => x"00",
  1481 => x"20",
  1482 => x"33",
  1483 => x"7c",
  1484 => x"00",
  1485 => x"ff",
  1486 => x"00",
  1487 => x"24",
  1488 => x"51",
  1489 => x"c9",
  1490 => x"ff",
  1491 => x"f8",
  1492 => x"34",
  1493 => x"3c",
  1494 => x"00",
  1495 => x"32",
  1496 => x"61",
  1497 => x"00",
  1498 => x"fe",
  1499 => x"96",
  1500 => x"3f",
  1501 => x"69",
  1502 => x"00",
  1503 => x"24",
  1504 => x"ff",
  1505 => x"fe",
  1506 => x"33",
  1507 => x"7c",
  1508 => x"00",
  1509 => x"00",
  1510 => x"00",
  1511 => x"22",
  1512 => x"b0",
  1513 => x"3c",
  1514 => x"00",
  1515 => x"01",
  1516 => x"67",
  1517 => x"12",
  1518 => x"51",
  1519 => x"ca",
  1520 => x"ff",
  1521 => x"e8",
  1522 => x"48",
  1523 => x"7a",
  1524 => x"ff",
  1525 => x"6e",
  1526 => x"61",
  1527 => x"00",
  1528 => x"01",
  1529 => x"22",
  1530 => x"58",
  1531 => x"8f",
  1532 => x"70",
  1533 => x"ff",
  1534 => x"4e",
  1535 => x"75",
  1536 => x"22",
  1537 => x"3c",
  1538 => x"00",
  1539 => x"00",
  1540 => x"20",
  1541 => x"00",
  1542 => x"33",
  1543 => x"7c",
  1544 => x"00",
  1545 => x"ff",
  1546 => x"00",
  1547 => x"24",
  1548 => x"53",
  1549 => x"81",
  1550 => x"66",
  1551 => x"f6",
  1552 => x"61",
  1553 => x"00",
  1554 => x"fe",
  1555 => x"72",
  1556 => x"b0",
  1557 => x"3c",
  1558 => x"00",
  1559 => x"01",
  1560 => x"66",
  1561 => x"00",
  1562 => x"00",
  1563 => x"9e",
  1564 => x"33",
  1565 => x"7c",
  1566 => x"00",
  1567 => x"ff",
  1568 => x"00",
  1569 => x"24",
  1570 => x"33",
  1571 => x"7c",
  1572 => x"00",
  1573 => x"ff",
  1574 => x"00",
  1575 => x"24",
  1576 => x"33",
  1577 => x"7c",
  1578 => x"00",
  1579 => x"ff",
  1580 => x"00",
  1581 => x"24",
  1582 => x"30",
  1583 => x"29",
  1584 => x"00",
  1585 => x"24",
  1586 => x"0c",
  1587 => x"00",
  1588 => x"00",
  1589 => x"01",
  1590 => x"66",
  1591 => x"00",
  1592 => x"00",
  1593 => x"80",
  1594 => x"33",
  1595 => x"7c",
  1596 => x"00",
  1597 => x"ff",
  1598 => x"00",
  1599 => x"24",
  1600 => x"30",
  1601 => x"29",
  1602 => x"00",
  1603 => x"24",
  1604 => x"0c",
  1605 => x"00",
  1606 => x"00",
  1607 => x"aa",
  1608 => x"66",
  1609 => x"6e",
  1610 => x"3f",
  1611 => x"69",
  1612 => x"00",
  1613 => x"24",
  1614 => x"ff",
  1615 => x"fe",
  1616 => x"33",
  1617 => x"7c",
  1618 => x"00",
  1619 => x"00",
  1620 => x"00",
  1621 => x"22",
  1622 => x"48",
  1623 => x"7a",
  1624 => x"ff",
  1625 => x"42",
  1626 => x"61",
  1627 => x"00",
  1628 => x"00",
  1629 => x"be",
  1630 => x"58",
  1631 => x"8f",
  1632 => x"34",
  1633 => x"3c",
  1634 => x"00",
  1635 => x"32",
  1636 => x"53",
  1637 => x"42",
  1638 => x"67",
  1639 => x"50",
  1640 => x"32",
  1641 => x"3c",
  1642 => x"07",
  1643 => x"d0",
  1644 => x"33",
  1645 => x"7c",
  1646 => x"00",
  1647 => x"ff",
  1648 => x"00",
  1649 => x"24",
  1650 => x"51",
  1651 => x"c9",
  1652 => x"ff",
  1653 => x"f8",
  1654 => x"61",
  1655 => x"00",
  1656 => x"fe",
  1657 => x"28",
  1658 => x"b0",
  1659 => x"3c",
  1660 => x"00",
  1661 => x"01",
  1662 => x"66",
  1663 => x"e4",
  1664 => x"61",
  1665 => x"00",
  1666 => x"fe",
  1667 => x"10",
  1668 => x"66",
  1669 => x"de",
  1670 => x"61",
  1671 => x"00",
  1672 => x"fe",
  1673 => x"22",
  1674 => x"66",
  1675 => x"d8",
  1676 => x"33",
  1677 => x"7c",
  1678 => x"00",
  1679 => x"ff",
  1680 => x"00",
  1681 => x"24",
  1682 => x"30",
  1683 => x"29",
  1684 => x"00",
  1685 => x"24",
  1686 => x"c0",
  1687 => x"3c",
  1688 => x"00",
  1689 => x"40",
  1690 => x"66",
  1691 => x"08",
  1692 => x"33",
  1693 => x"fc",
  1694 => x"00",
  1695 => x"00",
  1696 => x"00",
  1697 => x"7f",
  1698 => x"00",
  1699 => x"24",
  1700 => x"33",
  1701 => x"7c",
  1702 => x"00",
  1703 => x"ff",
  1704 => x"00",
  1705 => x"24",
  1706 => x"33",
  1707 => x"7c",
  1708 => x"00",
  1709 => x"ff",
  1710 => x"00",
  1711 => x"24",
  1712 => x"33",
  1713 => x"7c",
  1714 => x"00",
  1715 => x"ff",
  1716 => x"00",
  1717 => x"24",
  1718 => x"60",
  1719 => x"3c",
  1720 => x"33",
  1721 => x"fc",
  1722 => x"00",
  1723 => x"00",
  1724 => x"00",
  1725 => x"7f",
  1726 => x"00",
  1727 => x"24",
  1728 => x"34",
  1729 => x"3c",
  1730 => x"00",
  1731 => x"0a",
  1732 => x"32",
  1733 => x"3c",
  1734 => x"07",
  1735 => x"d0",
  1736 => x"33",
  1737 => x"7c",
  1738 => x"00",
  1739 => x"ff",
  1740 => x"00",
  1741 => x"24",
  1742 => x"51",
  1743 => x"c9",
  1744 => x"ff",
  1745 => x"f8",
  1746 => x"61",
  1747 => x"00",
  1748 => x"fd",
  1749 => x"a6",
  1750 => x"67",
  1751 => x"1c",
  1752 => x"3f",
  1753 => x"69",
  1754 => x"00",
  1755 => x"24",
  1756 => x"ff",
  1757 => x"fe",
  1758 => x"33",
  1759 => x"7c",
  1760 => x"00",
  1761 => x"00",
  1762 => x"00",
  1763 => x"22",
  1764 => x"51",
  1765 => x"ca",
  1766 => x"ff",
  1767 => x"de",
  1768 => x"48",
  1769 => x"7a",
  1770 => x"fe",
  1771 => x"69",
  1772 => x"61",
  1773 => x"2c",
  1774 => x"58",
  1775 => x"8f",
  1776 => x"70",
  1777 => x"ff",
  1778 => x"4e",
  1779 => x"75",
  1780 => x"3f",
  1781 => x"69",
  1782 => x"00",
  1783 => x"24",
  1784 => x"ff",
  1785 => x"fe",
  1786 => x"33",
  1787 => x"7c",
  1788 => x"00",
  1789 => x"00",
  1790 => x"00",
  1791 => x"22",
  1792 => x"33",
  1793 => x"69",
  1794 => x"00",
  1795 => x"2c",
  1796 => x"00",
  1797 => x"1e",
  1798 => x"48",
  1799 => x"7a",
  1800 => x"fe",
  1801 => x"3f",
  1802 => x"61",
  1803 => x"0e",
  1804 => x"58",
  1805 => x"8f",
  1806 => x"33",
  1807 => x"fc",
  1808 => x"ff",
  1809 => x"ff",
  1810 => x"81",
  1811 => x"00",
  1812 => x"00",
  1813 => x"06",
  1814 => x"70",
  1815 => x"00",
  1816 => x"4e",
  1817 => x"75",
  1818 => x"2f",
  1819 => x"08",
  1820 => x"20",
  1821 => x"6f",
  1822 => x"00",
  1823 => x"08",
  1824 => x"61",
  1825 => x"04",
  1826 => x"20",
  1827 => x"5f",
  1828 => x"4e",
  1829 => x"75",
  1830 => x"48",
  1831 => x"e7",
  1832 => x"00",
  1833 => x"c0",
  1834 => x"22",
  1835 => x"39",
  1836 => x"00",
  1837 => x"7f",
  1838 => x"00",
  1839 => x"52",
  1840 => x"43",
  1841 => x"f9",
  1842 => x"80",
  1843 => x"00",
  1844 => x"08",
  1845 => x"00",
  1846 => x"10",
  1847 => x"18",
  1848 => x"67",
  1849 => x"08",
  1850 => x"13",
  1851 => x"80",
  1852 => x"10",
  1853 => x"00",
  1854 => x"52",
  1855 => x"41",
  1856 => x"60",
  1857 => x"f4",
  1858 => x"06",
  1859 => x"b9",
  1860 => x"00",
  1861 => x"00",
  1862 => x"00",
  1863 => x"4c",
  1864 => x"00",
  1865 => x"7f",
  1866 => x"00",
  1867 => x"52",
  1868 => x"4c",
  1869 => x"df",
  1870 => x"03",
  1871 => x"00",
  1872 => x"4e",
  1873 => x"75",
  1874 => x"4a",
  1875 => x"79",
  1876 => x"00",
  1877 => x"7f",
  1878 => x"00",
  1879 => x"24",
  1880 => x"67",
  1881 => x"1e",
  1882 => x"41",
  1883 => x"fa",
  1884 => x"00",
  1885 => x"08",
  1886 => x"48",
  1887 => x"7a",
  1888 => x"00",
  1889 => x"34",
  1890 => x"60",
  1891 => x"c2",
  1892 => x"53",
  1893 => x"44",
  1894 => x"48",
  1895 => x"43",
  1896 => x"20",
  1897 => x"66",
  1898 => x"6c",
  1899 => x"61",
  1900 => x"67",
  1901 => x"20",
  1902 => x"73",
  1903 => x"74",
  1904 => x"69",
  1905 => x"6c",
  1906 => x"6c",
  1907 => x"20",
  1908 => x"73",
  1909 => x"65",
  1910 => x"74",
  1911 => x"00",
  1912 => x"41",
  1913 => x"fa",
  1914 => x"00",
  1915 => x"08",
  1916 => x"48",
  1917 => x"7a",
  1918 => x"00",
  1919 => x"16",
  1920 => x"60",
  1921 => x"a4",
  1922 => x"53",
  1923 => x"44",
  1924 => x"48",
  1925 => x"43",
  1926 => x"20",
  1927 => x"66",
  1928 => x"6c",
  1929 => x"61",
  1930 => x"67",
  1931 => x"20",
  1932 => x"63",
  1933 => x"6c",
  1934 => x"65",
  1935 => x"61",
  1936 => x"72",
  1937 => x"65",
  1938 => x"64",
  1939 => x"00",
  1940 => x"61",
  1941 => x"00",
  1942 => x"02",
  1943 => x"0a",
  1944 => x"61",
  1945 => x"00",
  1946 => x"fc",
  1947 => x"46",
  1948 => x"66",
  1949 => x"46",
  1950 => x"2e",
  1951 => x"3c",
  1952 => x"00",
  1953 => x"00",
  1954 => x"01",
  1955 => x"ff",
  1956 => x"41",
  1957 => x"f9",
  1958 => x"00",
  1959 => x"7f",
  1960 => x"00",
  1961 => x"56",
  1962 => x"43",
  1963 => x"f9",
  1964 => x"80",
  1965 => x"00",
  1966 => x"08",
  1967 => x"00",
  1968 => x"10",
  1969 => x"18",
  1970 => x"12",
  1971 => x"c0",
  1972 => x"48",
  1973 => x"e7",
  1974 => x"01",
  1975 => x"c0",
  1976 => x"61",
  1977 => x"00",
  1978 => x"f9",
  1979 => x"70",
  1980 => x"4c",
  1981 => x"df",
  1982 => x"03",
  1983 => x"80",
  1984 => x"51",
  1985 => x"cf",
  1986 => x"ff",
  1987 => x"ee",
  1988 => x"20",
  1989 => x"39",
  1990 => x"00",
  1991 => x"7f",
  1992 => x"00",
  1993 => x"38",
  1994 => x"52",
  1995 => x"80",
  1996 => x"23",
  1997 => x"c0",
  1998 => x"00",
  1999 => x"7f",
  2000 => x"00",
  2001 => x"38",
  2002 => x"53",
  2003 => x"79",
  2004 => x"00",
  2005 => x"7f",
  2006 => x"00",
  2007 => x"36",
  2008 => x"66",
  2009 => x"be",
  2010 => x"61",
  2011 => x"00",
  2012 => x"02",
  2013 => x"7a",
  2014 => x"66",
  2015 => x"b4",
  2016 => x"20",
  2017 => x"08",
  2018 => x"4e",
  2019 => x"75",
  2020 => x"70",
  2021 => x"00",
  2022 => x"4e",
  2023 => x"75",
  2024 => x"33",
  2025 => x"fc",
  2026 => x"02",
  2027 => x"01",
  2028 => x"81",
  2029 => x"00",
  2030 => x"00",
  2031 => x"06",
  2032 => x"70",
  2033 => x"00",
  2034 => x"23",
  2035 => x"c0",
  2036 => x"00",
  2037 => x"7f",
  2038 => x"00",
  2039 => x"3e",
  2040 => x"33",
  2041 => x"fc",
  2042 => x"02",
  2043 => x"11",
  2044 => x"81",
  2045 => x"00",
  2046 => x"00",
  2047 => x"06",
  2048 => x"61",
  2049 => x"00",
  2050 => x"fb",
  2051 => x"de",
  2052 => x"66",
  2053 => x"5c",
  2054 => x"33",
  2055 => x"fc",
  2056 => x"02",
  2057 => x"02",
  2058 => x"81",
  2059 => x"00",
  2060 => x"00",
  2061 => x"06",
  2062 => x"0c",
  2063 => x"28",
  2064 => x"00",
  2065 => x"55",
  2066 => x"01",
  2067 => x"fe",
  2068 => x"66",
  2069 => x"4c",
  2070 => x"0c",
  2071 => x"28",
  2072 => x"00",
  2073 => x"aa",
  2074 => x"01",
  2075 => x"ff",
  2076 => x"66",
  2077 => x"44",
  2078 => x"30",
  2079 => x"39",
  2080 => x"00",
  2081 => x"7f",
  2082 => x"00",
  2083 => x"26",
  2084 => x"c0",
  2085 => x"7c",
  2086 => x"00",
  2087 => x"70",
  2088 => x"b0",
  2089 => x"7c",
  2090 => x"00",
  2091 => x"40",
  2092 => x"64",
  2093 => x"40",
  2094 => x"43",
  2095 => x"e8",
  2096 => x"01",
  2097 => x"be",
  2098 => x"d2",
  2099 => x"c0",
  2100 => x"33",
  2101 => x"fc",
  2102 => x"02",
  2103 => x"03",
  2104 => x"81",
  2105 => x"00",
  2106 => x"00",
  2107 => x"06",
  2108 => x"20",
  2109 => x"29",
  2110 => x"00",
  2111 => x"08",
  2112 => x"e0",
  2113 => x"58",
  2114 => x"48",
  2115 => x"40",
  2116 => x"e0",
  2117 => x"58",
  2118 => x"23",
  2119 => x"c0",
  2120 => x"00",
  2121 => x"7f",
  2122 => x"00",
  2123 => x"3e",
  2124 => x"61",
  2125 => x"00",
  2126 => x"fb",
  2127 => x"92",
  2128 => x"66",
  2129 => x"10",
  2130 => x"0c",
  2131 => x"28",
  2132 => x"00",
  2133 => x"55",
  2134 => x"01",
  2135 => x"fe",
  2136 => x"66",
  2137 => x"08",
  2138 => x"0c",
  2139 => x"28",
  2140 => x"00",
  2141 => x"aa",
  2142 => x"01",
  2143 => x"ff",
  2144 => x"67",
  2145 => x"0c",
  2146 => x"33",
  2147 => x"fc",
  2148 => x"f2",
  2149 => x"01",
  2150 => x"81",
  2151 => x"00",
  2152 => x"00",
  2153 => x"06",
  2154 => x"70",
  2155 => x"ff",
  2156 => x"4e",
  2157 => x"75",
  2158 => x"33",
  2159 => x"fc",
  2160 => x"02",
  2161 => x"04",
  2162 => x"81",
  2163 => x"00",
  2164 => x"00",
  2165 => x"06",
  2166 => x"0c",
  2167 => x"a8",
  2168 => x"46",
  2169 => x"41",
  2170 => x"54",
  2171 => x"31",
  2172 => x"00",
  2173 => x"36",
  2174 => x"66",
  2175 => x"24",
  2176 => x"13",
  2177 => x"fc",
  2178 => x"00",
  2179 => x"0c",
  2180 => x"00",
  2181 => x"7f",
  2182 => x"00",
  2183 => x"28",
  2184 => x"0c",
  2185 => x"a8",
  2186 => x"32",
  2187 => x"20",
  2188 => x"20",
  2189 => x"20",
  2190 => x"00",
  2191 => x"3a",
  2192 => x"67",
  2193 => x"36",
  2194 => x"13",
  2195 => x"fc",
  2196 => x"00",
  2197 => x"10",
  2198 => x"00",
  2199 => x"7f",
  2200 => x"00",
  2201 => x"28",
  2202 => x"0c",
  2203 => x"a8",
  2204 => x"36",
  2205 => x"20",
  2206 => x"20",
  2207 => x"20",
  2208 => x"00",
  2209 => x"3a",
  2210 => x"67",
  2211 => x"24",
  2212 => x"13",
  2213 => x"fc",
  2214 => x"00",
  2215 => x"00",
  2216 => x"00",
  2217 => x"7f",
  2218 => x"00",
  2219 => x"28",
  2220 => x"0c",
  2221 => x"a8",
  2222 => x"46",
  2223 => x"41",
  2224 => x"54",
  2225 => x"33",
  2226 => x"00",
  2227 => x"52",
  2228 => x"66",
  2229 => x"ac",
  2230 => x"0c",
  2231 => x"a8",
  2232 => x"32",
  2233 => x"20",
  2234 => x"20",
  2235 => x"20",
  2236 => x"00",
  2237 => x"56",
  2238 => x"66",
  2239 => x"a2",
  2240 => x"13",
  2241 => x"fc",
  2242 => x"00",
  2243 => x"20",
  2244 => x"00",
  2245 => x"7f",
  2246 => x"00",
  2247 => x"28",
  2248 => x"20",
  2249 => x"28",
  2250 => x"00",
  2251 => x"0a",
  2252 => x"c0",
  2253 => x"bc",
  2254 => x"00",
  2255 => x"ff",
  2256 => x"ff",
  2257 => x"00",
  2258 => x"0c",
  2259 => x"80",
  2260 => x"00",
  2261 => x"00",
  2262 => x"02",
  2263 => x"00",
  2264 => x"66",
  2265 => x"88",
  2266 => x"22",
  2267 => x"39",
  2268 => x"00",
  2269 => x"7f",
  2270 => x"00",
  2271 => x"3e",
  2272 => x"30",
  2273 => x"28",
  2274 => x"00",
  2275 => x"0e",
  2276 => x"e0",
  2277 => x"58",
  2278 => x"d2",
  2279 => x"80",
  2280 => x"23",
  2281 => x"c1",
  2282 => x"00",
  2283 => x"7f",
  2284 => x"00",
  2285 => x"42",
  2286 => x"0c",
  2287 => x"39",
  2288 => x"00",
  2289 => x"20",
  2290 => x"00",
  2291 => x"7f",
  2292 => x"00",
  2293 => x"28",
  2294 => x"66",
  2295 => x"24",
  2296 => x"20",
  2297 => x"28",
  2298 => x"00",
  2299 => x"2c",
  2300 => x"e0",
  2301 => x"58",
  2302 => x"48",
  2303 => x"40",
  2304 => x"e0",
  2305 => x"58",
  2306 => x"23",
  2307 => x"c0",
  2308 => x"00",
  2309 => x"7f",
  2310 => x"00",
  2311 => x"2a",
  2312 => x"20",
  2313 => x"28",
  2314 => x"00",
  2315 => x"24",
  2316 => x"e0",
  2317 => x"58",
  2318 => x"48",
  2319 => x"40",
  2320 => x"e0",
  2321 => x"58",
  2322 => x"d2",
  2323 => x"80",
  2324 => x"53",
  2325 => x"28",
  2326 => x"00",
  2327 => x"10",
  2328 => x"66",
  2329 => x"f8",
  2330 => x"60",
  2331 => x"32",
  2332 => x"70",
  2333 => x"00",
  2334 => x"23",
  2335 => x"c0",
  2336 => x"00",
  2337 => x"7f",
  2338 => x"00",
  2339 => x"2a",
  2340 => x"30",
  2341 => x"28",
  2342 => x"00",
  2343 => x"16",
  2344 => x"e0",
  2345 => x"58",
  2346 => x"d2",
  2347 => x"80",
  2348 => x"53",
  2349 => x"28",
  2350 => x"00",
  2351 => x"10",
  2352 => x"66",
  2353 => x"f8",
  2354 => x"23",
  2355 => x"c1",
  2356 => x"00",
  2357 => x"7f",
  2358 => x"00",
  2359 => x"2e",
  2360 => x"20",
  2361 => x"01",
  2362 => x"10",
  2363 => x"28",
  2364 => x"00",
  2365 => x"12",
  2366 => x"e1",
  2367 => x"48",
  2368 => x"10",
  2369 => x"28",
  2370 => x"00",
  2371 => x"11",
  2372 => x"33",
  2373 => x"c0",
  2374 => x"00",
  2375 => x"7f",
  2376 => x"00",
  2377 => x"4e",
  2378 => x"e8",
  2379 => x"48",
  2380 => x"d2",
  2381 => x"80",
  2382 => x"70",
  2383 => x"00",
  2384 => x"10",
  2385 => x"28",
  2386 => x"00",
  2387 => x"0d",
  2388 => x"33",
  2389 => x"c0",
  2390 => x"00",
  2391 => x"7f",
  2392 => x"00",
  2393 => x"4a",
  2394 => x"92",
  2395 => x"80",
  2396 => x"92",
  2397 => x"80",
  2398 => x"23",
  2399 => x"c1",
  2400 => x"00",
  2401 => x"7f",
  2402 => x"00",
  2403 => x"46",
  2404 => x"33",
  2405 => x"fc",
  2406 => x"02",
  2407 => x"05",
  2408 => x"81",
  2409 => x"00",
  2410 => x"00",
  2411 => x"06",
  2412 => x"70",
  2413 => x"00",
  2414 => x"4e",
  2415 => x"75",
  2416 => x"20",
  2417 => x"39",
  2418 => x"00",
  2419 => x"7f",
  2420 => x"00",
  2421 => x"2a",
  2422 => x"23",
  2423 => x"c0",
  2424 => x"00",
  2425 => x"7f",
  2426 => x"00",
  2427 => x"32",
  2428 => x"66",
  2429 => x"28",
  2430 => x"42",
  2431 => x"b9",
  2432 => x"00",
  2433 => x"7f",
  2434 => x"00",
  2435 => x"32",
  2436 => x"30",
  2437 => x"39",
  2438 => x"00",
  2439 => x"7f",
  2440 => x"00",
  2441 => x"4e",
  2442 => x"e8",
  2443 => x"48",
  2444 => x"33",
  2445 => x"c0",
  2446 => x"00",
  2447 => x"7f",
  2448 => x"00",
  2449 => x"36",
  2450 => x"20",
  2451 => x"39",
  2452 => x"00",
  2453 => x"7f",
  2454 => x"00",
  2455 => x"2e",
  2456 => x"23",
  2457 => x"c0",
  2458 => x"00",
  2459 => x"7f",
  2460 => x"00",
  2461 => x"38",
  2462 => x"4e",
  2463 => x"75",
  2464 => x"20",
  2465 => x"39",
  2466 => x"00",
  2467 => x"7f",
  2468 => x"00",
  2469 => x"32",
  2470 => x"32",
  2471 => x"39",
  2472 => x"00",
  2473 => x"7f",
  2474 => x"00",
  2475 => x"4a",
  2476 => x"33",
  2477 => x"c1",
  2478 => x"00",
  2479 => x"7f",
  2480 => x"00",
  2481 => x"36",
  2482 => x"e2",
  2483 => x"49",
  2484 => x"65",
  2485 => x"04",
  2486 => x"e3",
  2487 => x"88",
  2488 => x"60",
  2489 => x"f8",
  2490 => x"d0",
  2491 => x"b9",
  2492 => x"00",
  2493 => x"7f",
  2494 => x"00",
  2495 => x"46",
  2496 => x"23",
  2497 => x"c0",
  2498 => x"00",
  2499 => x"7f",
  2500 => x"00",
  2501 => x"38",
  2502 => x"4e",
  2503 => x"75",
  2504 => x"48",
  2505 => x"e7",
  2506 => x"20",
  2507 => x"20",
  2508 => x"24",
  2509 => x"49",
  2510 => x"61",
  2511 => x"00",
  2512 => x"fa",
  2513 => x"10",
  2514 => x"66",
  2515 => x"7a",
  2516 => x"74",
  2517 => x"0f",
  2518 => x"4a",
  2519 => x"10",
  2520 => x"67",
  2521 => x"74",
  2522 => x"70",
  2523 => x"0a",
  2524 => x"12",
  2525 => x"32",
  2526 => x"00",
  2527 => x"00",
  2528 => x"b2",
  2529 => x"30",
  2530 => x"00",
  2531 => x"00",
  2532 => x"67",
  2533 => x"0a",
  2534 => x"d2",
  2535 => x"3c",
  2536 => x"00",
  2537 => x"20",
  2538 => x"b2",
  2539 => x"30",
  2540 => x"00",
  2541 => x"00",
  2542 => x"66",
  2543 => x"36",
  2544 => x"51",
  2545 => x"c8",
  2546 => x"ff",
  2547 => x"ea",
  2548 => x"70",
  2549 => x"00",
  2550 => x"10",
  2551 => x"28",
  2552 => x"00",
  2553 => x"0b",
  2554 => x"33",
  2555 => x"c0",
  2556 => x"00",
  2557 => x"7f",
  2558 => x"00",
  2559 => x"3c",
  2560 => x"0c",
  2561 => x"39",
  2562 => x"00",
  2563 => x"20",
  2564 => x"00",
  2565 => x"7f",
  2566 => x"00",
  2567 => x"28",
  2568 => x"66",
  2569 => x"08",
  2570 => x"30",
  2571 => x"28",
  2572 => x"00",
  2573 => x"14",
  2574 => x"e0",
  2575 => x"58",
  2576 => x"48",
  2577 => x"40",
  2578 => x"30",
  2579 => x"28",
  2580 => x"00",
  2581 => x"1a",
  2582 => x"e0",
  2583 => x"58",
  2584 => x"23",
  2585 => x"c0",
  2586 => x"00",
  2587 => x"7f",
  2588 => x"00",
  2589 => x"32",
  2590 => x"4c",
  2591 => x"df",
  2592 => x"04",
  2593 => x"04",
  2594 => x"70",
  2595 => x"ff",
  2596 => x"4e",
  2597 => x"75",
  2598 => x"41",
  2599 => x"e8",
  2600 => x"00",
  2601 => x"20",
  2602 => x"51",
  2603 => x"ca",
  2604 => x"ff",
  2605 => x"aa",
  2606 => x"20",
  2607 => x"39",
  2608 => x"00",
  2609 => x"7f",
  2610 => x"00",
  2611 => x"38",
  2612 => x"52",
  2613 => x"80",
  2614 => x"23",
  2615 => x"c0",
  2616 => x"00",
  2617 => x"7f",
  2618 => x"00",
  2619 => x"38",
  2620 => x"53",
  2621 => x"79",
  2622 => x"00",
  2623 => x"7f",
  2624 => x"00",
  2625 => x"36",
  2626 => x"66",
  2627 => x"8a",
  2628 => x"61",
  2629 => x"10",
  2630 => x"67",
  2631 => x"06",
  2632 => x"61",
  2633 => x"00",
  2634 => x"ff",
  2635 => x"56",
  2636 => x"60",
  2637 => x"80",
  2638 => x"4c",
  2639 => x"df",
  2640 => x"04",
  2641 => x"04",
  2642 => x"70",
  2643 => x"00",
  2644 => x"4e",
  2645 => x"75",
  2646 => x"0c",
  2647 => x"39",
  2648 => x"00",
  2649 => x"20",
  2650 => x"00",
  2651 => x"7f",
  2652 => x"00",
  2653 => x"28",
  2654 => x"67",
  2655 => x"3e",
  2656 => x"0c",
  2657 => x"39",
  2658 => x"00",
  2659 => x"0c",
  2660 => x"00",
  2661 => x"7f",
  2662 => x"00",
  2663 => x"28",
  2664 => x"67",
  2665 => x"78",
  2666 => x"20",
  2667 => x"39",
  2668 => x"00",
  2669 => x"7f",
  2670 => x"00",
  2671 => x"32",
  2672 => x"e0",
  2673 => x"88",
  2674 => x"d0",
  2675 => x"b9",
  2676 => x"00",
  2677 => x"7f",
  2678 => x"00",
  2679 => x"42",
  2680 => x"61",
  2681 => x"00",
  2682 => x"f9",
  2683 => x"66",
  2684 => x"66",
  2685 => x"60",
  2686 => x"10",
  2687 => x"39",
  2688 => x"00",
  2689 => x"7f",
  2690 => x"00",
  2691 => x"35",
  2692 => x"d0",
  2693 => x"40",
  2694 => x"30",
  2695 => x"30",
  2696 => x"00",
  2697 => x"00",
  2698 => x"e0",
  2699 => x"58",
  2700 => x"23",
  2701 => x"c0",
  2702 => x"00",
  2703 => x"7f",
  2704 => x"00",
  2705 => x"32",
  2706 => x"80",
  2707 => x"bc",
  2708 => x"ff",
  2709 => x"ff",
  2710 => x"00",
  2711 => x"0f",
  2712 => x"b0",
  2713 => x"7c",
  2714 => x"ff",
  2715 => x"ff",
  2716 => x"4e",
  2717 => x"75",
  2718 => x"20",
  2719 => x"39",
  2720 => x"00",
  2721 => x"7f",
  2722 => x"00",
  2723 => x"32",
  2724 => x"ee",
  2725 => x"88",
  2726 => x"d0",
  2727 => x"b9",
  2728 => x"00",
  2729 => x"7f",
  2730 => x"00",
  2731 => x"42",
  2732 => x"61",
  2733 => x"00",
  2734 => x"f9",
  2735 => x"32",
  2736 => x"66",
  2737 => x"2c",
  2738 => x"10",
  2739 => x"39",
  2740 => x"00",
  2741 => x"7f",
  2742 => x"00",
  2743 => x"35",
  2744 => x"c0",
  2745 => x"7c",
  2746 => x"00",
  2747 => x"7f",
  2748 => x"d0",
  2749 => x"40",
  2750 => x"d0",
  2751 => x"40",
  2752 => x"20",
  2753 => x"30",
  2754 => x"00",
  2755 => x"00",
  2756 => x"e0",
  2757 => x"58",
  2758 => x"48",
  2759 => x"40",
  2760 => x"e0",
  2761 => x"58",
  2762 => x"23",
  2763 => x"c0",
  2764 => x"00",
  2765 => x"7f",
  2766 => x"00",
  2767 => x"32",
  2768 => x"80",
  2769 => x"bc",
  2770 => x"f0",
  2771 => x"00",
  2772 => x"00",
  2773 => x"07",
  2774 => x"b0",
  2775 => x"bc",
  2776 => x"ff",
  2777 => x"ff",
  2778 => x"ff",
  2779 => x"ff",
  2780 => x"4e",
  2781 => x"75",
  2782 => x"70",
  2783 => x"00",
  2784 => x"4e",
  2785 => x"75",
  2786 => x"2f",
  2787 => x"02",
  2788 => x"20",
  2789 => x"39",
  2790 => x"00",
  2791 => x"7f",
  2792 => x"00",
  2793 => x"32",
  2794 => x"22",
  2795 => x"00",
  2796 => x"d0",
  2797 => x"80",
  2798 => x"d0",
  2799 => x"81",
  2800 => x"22",
  2801 => x"00",
  2802 => x"e0",
  2803 => x"88",
  2804 => x"e4",
  2805 => x"88",
  2806 => x"d0",
  2807 => x"b9",
  2808 => x"00",
  2809 => x"7f",
  2810 => x"00",
  2811 => x"42",
  2812 => x"24",
  2813 => x"00",
  2814 => x"61",
  2815 => x"00",
  2816 => x"f8",
  2817 => x"e0",
  2818 => x"66",
  2819 => x"52",
  2820 => x"20",
  2821 => x"01",
  2822 => x"e2",
  2823 => x"88",
  2824 => x"c0",
  2825 => x"7c",
  2826 => x"01",
  2827 => x"ff",
  2828 => x"b0",
  2829 => x"7c",
  2830 => x"01",
  2831 => x"ff",
  2832 => x"66",
  2833 => x"14",
  2834 => x"10",
  2835 => x"30",
  2836 => x"00",
  2837 => x"00",
  2838 => x"c1",
  2839 => x"42",
  2840 => x"52",
  2841 => x"80",
  2842 => x"61",
  2843 => x"00",
  2844 => x"f8",
  2845 => x"c4",
  2846 => x"66",
  2847 => x"36",
  2848 => x"e1",
  2849 => x"4a",
  2850 => x"14",
  2851 => x"10",
  2852 => x"60",
  2853 => x"0a",
  2854 => x"14",
  2855 => x"30",
  2856 => x"00",
  2857 => x"00",
  2858 => x"e1",
  2859 => x"4a",
  2860 => x"14",
  2861 => x"30",
  2862 => x"00",
  2863 => x"01",
  2864 => x"e1",
  2865 => x"5a",
  2866 => x"c2",
  2867 => x"7c",
  2868 => x"00",
  2869 => x"01",
  2870 => x"67",
  2871 => x"02",
  2872 => x"e8",
  2873 => x"4a",
  2874 => x"c4",
  2875 => x"bc",
  2876 => x"00",
  2877 => x"00",
  2878 => x"0f",
  2879 => x"ff",
  2880 => x"23",
  2881 => x"c2",
  2882 => x"00",
  2883 => x"7f",
  2884 => x"00",
  2885 => x"32",
  2886 => x"84",
  2887 => x"bc",
  2888 => x"ff",
  2889 => x"ff",
  2890 => x"f0",
  2891 => x"0f",
  2892 => x"20",
  2893 => x"02",
  2894 => x"24",
  2895 => x"1f",
  2896 => x"b0",
  2897 => x"7c",
  2898 => x"ff",
  2899 => x"ff",
  2900 => x"4e",
  2901 => x"75",
  2902 => x"24",
  2903 => x"1f",
  2904 => x"70",
  2905 => x"00",
  2906 => x"4e",
  2907 => x"75",
  2908 => x"41",
  2909 => x"f9",
  2910 => x"00",
  2911 => x"7f",
  2912 => x"00",
  2913 => x"04",
  2914 => x"20",
  2915 => x"bc",
  2916 => x"12",
  2917 => x"34",
  2918 => x"56",
  2919 => x"78",
  2920 => x"21",
  2921 => x"7c",
  2922 => x"fe",
  2923 => x"dc",
  2924 => x"ba",
  2925 => x"98",
  2926 => x"00",
  2927 => x"04",
  2928 => x"21",
  2929 => x"7c",
  2930 => x"aa",
  2931 => x"55",
  2932 => x"cc",
  2933 => x"22",
  2934 => x"00",
  2935 => x"02",
  2936 => x"11",
  2937 => x"7c",
  2938 => x"00",
  2939 => x"33",
  2940 => x"00",
  2941 => x"03",
  2942 => x"11",
  2943 => x"7c",
  2944 => x"00",
  2945 => x"fe",
  2946 => x"00",
  2947 => x"04",
  2948 => x"20",
  2949 => x"10",
  2950 => x"22",
  2951 => x"28",
  2952 => x"00",
  2953 => x"04",
  2954 => x"90",
  2955 => x"bc",
  2956 => x"12",
  2957 => x"34",
  2958 => x"aa",
  2959 => x"33",
  2960 => x"92",
  2961 => x"bc",
  2962 => x"fe",
  2963 => x"22",
  2964 => x"ba",
  2965 => x"98",
  2966 => x"80",
  2967 => x"81",
  2968 => x"4e",
  2969 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;


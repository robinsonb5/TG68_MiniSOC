library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Hex_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end Hex_ROM;

architecture arch of Hex_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"00",
     2 => x"0f",
     3 => x"fe",
     4 => x"00",
     5 => x"00",
     6 => x"01",
     7 => x"00",
     8 => x"00",
     9 => x"00",
    10 => x"00",
    11 => x"00",
    12 => x"00",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"00",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"00",
    21 => x"00",
    22 => x"00",
    23 => x"00",
    24 => x"00",
    25 => x"00",
    26 => x"00",
    27 => x"00",
    28 => x"00",
    29 => x"00",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"00",
    34 => x"00",
    35 => x"00",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"00",
    40 => x"00",
    41 => x"00",
    42 => x"00",
    43 => x"00",
    44 => x"00",
    45 => x"00",
    46 => x"00",
    47 => x"00",
    48 => x"00",
    49 => x"00",
    50 => x"00",
    51 => x"00",
    52 => x"00",
    53 => x"00",
    54 => x"00",
    55 => x"00",
    56 => x"00",
    57 => x"00",
    58 => x"00",
    59 => x"00",
    60 => x"00",
    61 => x"00",
    62 => x"00",
    63 => x"00",
    64 => x"00",
    65 => x"00",
    66 => x"00",
    67 => x"00",
    68 => x"00",
    69 => x"00",
    70 => x"00",
    71 => x"00",
    72 => x"00",
    73 => x"00",
    74 => x"00",
    75 => x"00",
    76 => x"00",
    77 => x"00",
    78 => x"00",
    79 => x"00",
    80 => x"00",
    81 => x"00",
    82 => x"00",
    83 => x"00",
    84 => x"00",
    85 => x"00",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"00",
    93 => x"00",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"00",
   127 => x"00",
   128 => x"00",
   129 => x"00",
   130 => x"00",
   131 => x"00",
   132 => x"00",
   133 => x"00",
   134 => x"00",
   135 => x"00",
   136 => x"00",
   137 => x"00",
   138 => x"00",
   139 => x"00",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"00",
   144 => x"00",
   145 => x"00",
   146 => x"00",
   147 => x"00",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"00",
   153 => x"00",
   154 => x"00",
   155 => x"00",
   156 => x"00",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"00",
   161 => x"00",
   162 => x"00",
   163 => x"00",
   164 => x"00",
   165 => x"00",
   166 => x"00",
   167 => x"00",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"00",
   172 => x"00",
   173 => x"00",
   174 => x"00",
   175 => x"00",
   176 => x"00",
   177 => x"00",
   178 => x"00",
   179 => x"00",
   180 => x"00",
   181 => x"00",
   182 => x"00",
   183 => x"00",
   184 => x"00",
   185 => x"00",
   186 => x"00",
   187 => x"00",
   188 => x"00",
   189 => x"00",
   190 => x"00",
   191 => x"00",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"00",
   196 => x"00",
   197 => x"00",
   198 => x"00",
   199 => x"00",
   200 => x"00",
   201 => x"00",
   202 => x"00",
   203 => x"00",
   204 => x"00",
   205 => x"00",
   206 => x"00",
   207 => x"00",
   208 => x"00",
   209 => x"00",
   210 => x"00",
   211 => x"00",
   212 => x"00",
   213 => x"00",
   214 => x"00",
   215 => x"00",
   216 => x"00",
   217 => x"00",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"00",
   224 => x"00",
   225 => x"00",
   226 => x"00",
   227 => x"00",
   228 => x"00",
   229 => x"00",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"00",
   234 => x"00",
   235 => x"00",
   236 => x"00",
   237 => x"00",
   238 => x"00",
   239 => x"00",
   240 => x"00",
   241 => x"00",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"00",
   248 => x"00",
   249 => x"00",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"00",
   256 => x"4f",
   257 => x"f9",
   258 => x"00",
   259 => x"00",
   260 => x"0f",
   261 => x"fe",
   262 => x"41",
   263 => x"f9",
   264 => x"00",
   265 => x"00",
   266 => x"0c",
   267 => x"48",
   268 => x"20",
   269 => x"3c",
   270 => x"00",
   271 => x"00",
   272 => x"0c",
   273 => x"48",
   274 => x"b1",
   275 => x"c0",
   276 => x"6c",
   277 => x"04",
   278 => x"42",
   279 => x"98",
   280 => x"60",
   281 => x"f8",
   282 => x"41",
   283 => x"fa",
   284 => x"00",
   285 => x"4e",
   286 => x"21",
   287 => x"c8",
   288 => x"00",
   289 => x"64",
   290 => x"41",
   291 => x"fa",
   292 => x"00",
   293 => x"54",
   294 => x"21",
   295 => x"c8",
   296 => x"00",
   297 => x"68",
   298 => x"41",
   299 => x"fa",
   300 => x"00",
   301 => x"5a",
   302 => x"21",
   303 => x"c8",
   304 => x"00",
   305 => x"6c",
   306 => x"41",
   307 => x"fa",
   308 => x"00",
   309 => x"60",
   310 => x"21",
   311 => x"c8",
   312 => x"00",
   313 => x"70",
   314 => x"41",
   315 => x"fa",
   316 => x"00",
   317 => x"66",
   318 => x"21",
   319 => x"c8",
   320 => x"00",
   321 => x"74",
   322 => x"41",
   323 => x"fa",
   324 => x"00",
   325 => x"6c",
   326 => x"21",
   327 => x"c8",
   328 => x"00",
   329 => x"78",
   330 => x"41",
   331 => x"fa",
   332 => x"00",
   333 => x"72",
   334 => x"21",
   335 => x"c8",
   336 => x"00",
   337 => x"7c",
   338 => x"48",
   339 => x"78",
   340 => x"00",
   341 => x"01",
   342 => x"48",
   343 => x"7a",
   344 => x"00",
   345 => x"0a",
   346 => x"4e",
   347 => x"b9",
   348 => x"00",
   349 => x"00",
   350 => x"02",
   351 => x"80",
   352 => x"60",
   353 => x"fe",
   354 => x"42",
   355 => x"6f",
   356 => x"6f",
   357 => x"74",
   358 => x"72",
   359 => x"6f",
   360 => x"6d",
   361 => x"00",
   362 => x"48",
   363 => x"e7",
   364 => x"ff",
   365 => x"fe",
   366 => x"48",
   367 => x"7a",
   368 => x"00",
   369 => x"5c",
   370 => x"2f",
   371 => x"3a",
   372 => x"00",
   373 => x"60",
   374 => x"4e",
   375 => x"75",
   376 => x"48",
   377 => x"e7",
   378 => x"ff",
   379 => x"fe",
   380 => x"48",
   381 => x"7a",
   382 => x"00",
   383 => x"4e",
   384 => x"2f",
   385 => x"3a",
   386 => x"00",
   387 => x"56",
   388 => x"4e",
   389 => x"75",
   390 => x"48",
   391 => x"e7",
   392 => x"ff",
   393 => x"fe",
   394 => x"48",
   395 => x"7a",
   396 => x"00",
   397 => x"40",
   398 => x"2f",
   399 => x"3a",
   400 => x"00",
   401 => x"4c",
   402 => x"4e",
   403 => x"75",
   404 => x"48",
   405 => x"e7",
   406 => x"ff",
   407 => x"fe",
   408 => x"48",
   409 => x"7a",
   410 => x"00",
   411 => x"32",
   412 => x"2f",
   413 => x"3a",
   414 => x"00",
   415 => x"42",
   416 => x"4e",
   417 => x"75",
   418 => x"48",
   419 => x"e7",
   420 => x"ff",
   421 => x"fe",
   422 => x"48",
   423 => x"7a",
   424 => x"00",
   425 => x"24",
   426 => x"2f",
   427 => x"3a",
   428 => x"00",
   429 => x"38",
   430 => x"4e",
   431 => x"75",
   432 => x"48",
   433 => x"e7",
   434 => x"ff",
   435 => x"fe",
   436 => x"48",
   437 => x"7a",
   438 => x"00",
   439 => x"16",
   440 => x"2f",
   441 => x"3a",
   442 => x"00",
   443 => x"2e",
   444 => x"4e",
   445 => x"75",
   446 => x"48",
   447 => x"e7",
   448 => x"ff",
   449 => x"fe",
   450 => x"48",
   451 => x"7a",
   452 => x"00",
   453 => x"08",
   454 => x"2f",
   455 => x"3a",
   456 => x"00",
   457 => x"24",
   458 => x"4e",
   459 => x"75",
   460 => x"4c",
   461 => x"df",
   462 => x"7f",
   463 => x"ff",
   464 => x"4e",
   465 => x"73",
   466 => x"4e",
   467 => x"75",
   468 => x"00",
   469 => x"00",
   470 => x"01",
   471 => x"d2",
   472 => x"00",
   473 => x"00",
   474 => x"01",
   475 => x"d2",
   476 => x"00",
   477 => x"00",
   478 => x"01",
   479 => x"d2",
   480 => x"00",
   481 => x"00",
   482 => x"01",
   483 => x"d2",
   484 => x"00",
   485 => x"00",
   486 => x"01",
   487 => x"d2",
   488 => x"00",
   489 => x"00",
   490 => x"01",
   491 => x"d2",
   492 => x"00",
   493 => x"00",
   494 => x"01",
   495 => x"d2",
   496 => x"46",
   497 => x"fc",
   498 => x"20",
   499 => x"00",
   500 => x"4e",
   501 => x"75",
   502 => x"46",
   503 => x"fc",
   504 => x"27",
   505 => x"00",
   506 => x"4e",
   507 => x"75",
   508 => x"00",
   509 => x"00",
   510 => x"00",
   511 => x"00",
   512 => x"cf",
   513 => x"00",
   514 => x"00",
   515 => x"00",
   516 => x"00",
   517 => x"00",
   518 => x"00",
   519 => x"00",
   520 => x"8c",
   521 => x"ff",
   522 => x"f0",
   523 => x"00",
   524 => x"00",
   525 => x"00",
   526 => x"00",
   527 => x"00",
   528 => x"08",
   529 => x"cc",
   530 => x"ff",
   531 => x"f0",
   532 => x"00",
   533 => x"00",
   534 => x"00",
   535 => x"00",
   536 => x"08",
   537 => x"cc",
   538 => x"cc",
   539 => x"ff",
   540 => x"ff",
   541 => x"00",
   542 => x"00",
   543 => x"00",
   544 => x"08",
   545 => x"8c",
   546 => x"cc",
   547 => x"cc",
   548 => x"cf",
   549 => x"ff",
   550 => x"00",
   551 => x"00",
   552 => x"00",
   553 => x"8c",
   554 => x"cc",
   555 => x"cc",
   556 => x"cc",
   557 => x"c8",
   558 => x"00",
   559 => x"00",
   560 => x"00",
   561 => x"88",
   562 => x"cc",
   563 => x"cc",
   564 => x"cc",
   565 => x"80",
   566 => x"00",
   567 => x"00",
   568 => x"00",
   569 => x"08",
   570 => x"cc",
   571 => x"cc",
   572 => x"cf",
   573 => x"00",
   574 => x"00",
   575 => x"00",
   576 => x"00",
   577 => x"08",
   578 => x"cc",
   579 => x"cc",
   580 => x"cc",
   581 => x"f0",
   582 => x"00",
   583 => x"00",
   584 => x"00",
   585 => x"08",
   586 => x"8c",
   587 => x"c8",
   588 => x"cc",
   589 => x"cf",
   590 => x"00",
   591 => x"00",
   592 => x"00",
   593 => x"00",
   594 => x"8c",
   595 => x"80",
   596 => x"8c",
   597 => x"cc",
   598 => x"f0",
   599 => x"00",
   600 => x"00",
   601 => x"00",
   602 => x"88",
   603 => x"00",
   604 => x"08",
   605 => x"cc",
   606 => x"cf",
   607 => x"00",
   608 => x"00",
   609 => x"00",
   610 => x"00",
   611 => x"00",
   612 => x"00",
   613 => x"8c",
   614 => x"cc",
   615 => x"f0",
   616 => x"00",
   617 => x"00",
   618 => x"00",
   619 => x"00",
   620 => x"00",
   621 => x"08",
   622 => x"cc",
   623 => x"c8",
   624 => x"00",
   625 => x"00",
   626 => x"00",
   627 => x"00",
   628 => x"00",
   629 => x"00",
   630 => x"8c",
   631 => x"80",
   632 => x"00",
   633 => x"00",
   634 => x"00",
   635 => x"00",
   636 => x"00",
   637 => x"00",
   638 => x"08",
   639 => x"00",
   640 => x"4e",
   641 => x"56",
   642 => x"00",
   643 => x"00",
   644 => x"2f",
   645 => x"0a",
   646 => x"30",
   647 => x"39",
   648 => x"81",
   649 => x"00",
   650 => x"00",
   651 => x"2a",
   652 => x"48",
   653 => x"78",
   654 => x"04",
   655 => x"80",
   656 => x"c0",
   657 => x"fc",
   658 => x"03",
   659 => x"e8",
   660 => x"2f",
   661 => x"00",
   662 => x"4e",
   663 => x"b9",
   664 => x"00",
   665 => x"00",
   666 => x"08",
   667 => x"f8",
   668 => x"50",
   669 => x"8f",
   670 => x"33",
   671 => x"c0",
   672 => x"81",
   673 => x"00",
   674 => x"00",
   675 => x"02",
   676 => x"48",
   677 => x"79",
   678 => x"00",
   679 => x"00",
   680 => x"0b",
   681 => x"f2",
   682 => x"45",
   683 => x"f9",
   684 => x"00",
   685 => x"00",
   686 => x"03",
   687 => x"0e",
   688 => x"4e",
   689 => x"92",
   690 => x"48",
   691 => x"79",
   692 => x"00",
   693 => x"00",
   694 => x"0c",
   695 => x"00",
   696 => x"4e",
   697 => x"92",
   698 => x"2f",
   699 => x"3c",
   700 => x"00",
   701 => x"01",
   702 => x"00",
   703 => x"00",
   704 => x"4e",
   705 => x"b9",
   706 => x"00",
   707 => x"00",
   708 => x"07",
   709 => x"64",
   710 => x"4f",
   711 => x"ef",
   712 => x"00",
   713 => x"0c",
   714 => x"4a",
   715 => x"80",
   716 => x"67",
   717 => x"0e",
   718 => x"48",
   719 => x"79",
   720 => x"00",
   721 => x"00",
   722 => x"0c",
   723 => x"1d",
   724 => x"4e",
   725 => x"92",
   726 => x"58",
   727 => x"8f",
   728 => x"70",
   729 => x"00",
   730 => x"60",
   731 => x"08",
   732 => x"48",
   733 => x"79",
   734 => x"00",
   735 => x"00",
   736 => x"0c",
   737 => x"32",
   738 => x"60",
   739 => x"f0",
   740 => x"33",
   741 => x"c0",
   742 => x"81",
   743 => x"00",
   744 => x"00",
   745 => x"06",
   746 => x"52",
   747 => x"80",
   748 => x"60",
   749 => x"f6",
   750 => x"00",
   751 => x"00",
   752 => x"4e",
   753 => x"56",
   754 => x"00",
   755 => x"00",
   756 => x"20",
   757 => x"2e",
   758 => x"00",
   759 => x"08",
   760 => x"32",
   761 => x"39",
   762 => x"81",
   763 => x"00",
   764 => x"00",
   765 => x"00",
   766 => x"08",
   767 => x"01",
   768 => x"00",
   769 => x"08",
   770 => x"67",
   771 => x"f4",
   772 => x"33",
   773 => x"c0",
   774 => x"81",
   775 => x"00",
   776 => x"00",
   777 => x"00",
   778 => x"4e",
   779 => x"5e",
   780 => x"4e",
   781 => x"75",
   782 => x"4e",
   783 => x"56",
   784 => x"00",
   785 => x"00",
   786 => x"48",
   787 => x"e7",
   788 => x"20",
   789 => x"30",
   790 => x"24",
   791 => x"6e",
   792 => x"00",
   793 => x"08",
   794 => x"47",
   795 => x"fa",
   796 => x"ff",
   797 => x"d4",
   798 => x"60",
   799 => x"0c",
   800 => x"48",
   801 => x"80",
   802 => x"30",
   803 => x"40",
   804 => x"2f",
   805 => x"08",
   806 => x"4e",
   807 => x"93",
   808 => x"52",
   809 => x"82",
   810 => x"58",
   811 => x"8f",
   812 => x"10",
   813 => x"1a",
   814 => x"66",
   815 => x"f0",
   816 => x"20",
   817 => x"02",
   818 => x"4c",
   819 => x"ee",
   820 => x"0c",
   821 => x"04",
   822 => x"ff",
   823 => x"f4",
   824 => x"4e",
   825 => x"5e",
   826 => x"4e",
   827 => x"75",
   828 => x"4e",
   829 => x"56",
   830 => x"00",
   831 => x"00",
   832 => x"70",
   833 => x"00",
   834 => x"60",
   835 => x"0c",
   836 => x"30",
   837 => x"39",
   838 => x"81",
   839 => x"00",
   840 => x"00",
   841 => x"00",
   842 => x"02",
   843 => x"80",
   844 => x"00",
   845 => x"00",
   846 => x"ff",
   847 => x"ff",
   848 => x"08",
   849 => x"00",
   850 => x"00",
   851 => x"09",
   852 => x"67",
   853 => x"ee",
   854 => x"4e",
   855 => x"5e",
   856 => x"4e",
   857 => x"75",
   858 => x"00",
   859 => x"00",
   860 => x"4e",
   861 => x"56",
   862 => x"00",
   863 => x"00",
   864 => x"48",
   865 => x"e7",
   866 => x"38",
   867 => x"20",
   868 => x"24",
   869 => x"2e",
   870 => x"00",
   871 => x"08",
   872 => x"67",
   873 => x"3a",
   874 => x"76",
   875 => x"08",
   876 => x"70",
   877 => x"00",
   878 => x"45",
   879 => x"f9",
   880 => x"00",
   881 => x"00",
   882 => x"02",
   883 => x"f0",
   884 => x"22",
   885 => x"02",
   886 => x"78",
   887 => x"1c",
   888 => x"e8",
   889 => x"a9",
   890 => x"20",
   891 => x"41",
   892 => x"e9",
   893 => x"8a",
   894 => x"4a",
   895 => x"81",
   896 => x"67",
   897 => x"0c",
   898 => x"70",
   899 => x"09",
   900 => x"b0",
   901 => x"81",
   902 => x"6c",
   903 => x"0a",
   904 => x"41",
   905 => x"e8",
   906 => x"00",
   907 => x"37",
   908 => x"60",
   909 => x"08",
   910 => x"4a",
   911 => x"80",
   912 => x"67",
   913 => x"0c",
   914 => x"41",
   915 => x"e8",
   916 => x"00",
   917 => x"30",
   918 => x"2f",
   919 => x"08",
   920 => x"4e",
   921 => x"92",
   922 => x"58",
   923 => x"8f",
   924 => x"70",
   925 => x"01",
   926 => x"53",
   927 => x"83",
   928 => x"66",
   929 => x"d2",
   930 => x"60",
   931 => x"0c",
   932 => x"48",
   933 => x"78",
   934 => x"00",
   935 => x"30",
   936 => x"4e",
   937 => x"b9",
   938 => x"00",
   939 => x"00",
   940 => x"02",
   941 => x"f0",
   942 => x"58",
   943 => x"8f",
   944 => x"48",
   945 => x"78",
   946 => x"00",
   947 => x"0a",
   948 => x"4e",
   949 => x"b9",
   950 => x"00",
   951 => x"00",
   952 => x"02",
   953 => x"f0",
   954 => x"70",
   955 => x"00",
   956 => x"4c",
   957 => x"ee",
   958 => x"04",
   959 => x"1c",
   960 => x"ff",
   961 => x"f0",
   962 => x"4e",
   963 => x"5e",
   964 => x"4e",
   965 => x"75",
   966 => x"4e",
   967 => x"56",
   968 => x"00",
   969 => x"00",
   970 => x"20",
   971 => x"6e",
   972 => x"00",
   973 => x"08",
   974 => x"20",
   975 => x"28",
   976 => x"40",
   977 => x"00",
   978 => x"20",
   979 => x"3c",
   980 => x"00",
   981 => x"01",
   982 => x"00",
   983 => x"04",
   984 => x"20",
   985 => x"30",
   986 => x"08",
   987 => x"00",
   988 => x"20",
   989 => x"3c",
   990 => x"00",
   991 => x"00",
   992 => x"80",
   993 => x"00",
   994 => x"20",
   995 => x"30",
   996 => x"08",
   997 => x"00",
   998 => x"20",
   999 => x"3c",
  1000 => x"00",
  1001 => x"00",
  1002 => x"c0",
  1003 => x"0c",
  1004 => x"20",
  1005 => x"30",
  1006 => x"08",
  1007 => x"00",
  1008 => x"20",
  1009 => x"3c",
  1010 => x"00",
  1011 => x"00",
  1012 => x"c0",
  1013 => x"04",
  1014 => x"20",
  1015 => x"30",
  1016 => x"08",
  1017 => x"00",
  1018 => x"20",
  1019 => x"3c",
  1020 => x"00",
  1021 => x"00",
  1022 => x"80",
  1023 => x"0c",
  1024 => x"20",
  1025 => x"30",
  1026 => x"08",
  1027 => x"00",
  1028 => x"70",
  1029 => x"01",
  1030 => x"48",
  1031 => x"40",
  1032 => x"20",
  1033 => x"30",
  1034 => x"08",
  1035 => x"00",
  1036 => x"20",
  1037 => x"28",
  1038 => x"40",
  1039 => x"08",
  1040 => x"4e",
  1041 => x"5e",
  1042 => x"4e",
  1043 => x"75",
  1044 => x"4e",
  1045 => x"56",
  1046 => x"00",
  1047 => x"00",
  1048 => x"48",
  1049 => x"e7",
  1050 => x"38",
  1051 => x"20",
  1052 => x"24",
  1053 => x"6e",
  1054 => x"00",
  1055 => x"08",
  1056 => x"20",
  1057 => x"2e",
  1058 => x"00",
  1059 => x"0c",
  1060 => x"24",
  1061 => x"00",
  1062 => x"48",
  1063 => x"42",
  1064 => x"42",
  1065 => x"42",
  1066 => x"84",
  1067 => x"6e",
  1068 => x"00",
  1069 => x"10",
  1070 => x"24",
  1071 => x"80",
  1072 => x"25",
  1073 => x"6e",
  1074 => x"00",
  1075 => x"10",
  1076 => x"00",
  1077 => x"04",
  1078 => x"26",
  1079 => x"2a",
  1080 => x"00",
  1081 => x"02",
  1082 => x"b4",
  1083 => x"83",
  1084 => x"67",
  1085 => x"18",
  1086 => x"48",
  1087 => x"79",
  1088 => x"00",
  1089 => x"00",
  1090 => x"09",
  1091 => x"84",
  1092 => x"4e",
  1093 => x"b9",
  1094 => x"00",
  1095 => x"00",
  1096 => x"03",
  1097 => x"0e",
  1098 => x"2f",
  1099 => x"03",
  1100 => x"4e",
  1101 => x"ba",
  1102 => x"ff",
  1103 => x"0e",
  1104 => x"b5",
  1105 => x"83",
  1106 => x"50",
  1107 => x"8f",
  1108 => x"60",
  1109 => x"02",
  1110 => x"76",
  1111 => x"00",
  1112 => x"48",
  1113 => x"6a",
  1114 => x"00",
  1115 => x"08",
  1116 => x"4e",
  1117 => x"ba",
  1118 => x"ff",
  1119 => x"68",
  1120 => x"28",
  1121 => x"2a",
  1122 => x"00",
  1123 => x"02",
  1124 => x"58",
  1125 => x"8f",
  1126 => x"b4",
  1127 => x"84",
  1128 => x"67",
  1129 => x"18",
  1130 => x"48",
  1131 => x"79",
  1132 => x"00",
  1133 => x"00",
  1134 => x"09",
  1135 => x"ab",
  1136 => x"4e",
  1137 => x"b9",
  1138 => x"00",
  1139 => x"00",
  1140 => x"03",
  1141 => x"0e",
  1142 => x"2f",
  1143 => x"04",
  1144 => x"4e",
  1145 => x"ba",
  1146 => x"fe",
  1147 => x"e2",
  1148 => x"b9",
  1149 => x"82",
  1150 => x"86",
  1151 => x"82",
  1152 => x"50",
  1153 => x"8f",
  1154 => x"20",
  1155 => x"03",
  1156 => x"4c",
  1157 => x"ee",
  1158 => x"04",
  1159 => x"1c",
  1160 => x"ff",
  1161 => x"f0",
  1162 => x"4e",
  1163 => x"5e",
  1164 => x"4e",
  1165 => x"75",
  1166 => x"4e",
  1167 => x"56",
  1168 => x"00",
  1169 => x"00",
  1170 => x"48",
  1171 => x"e7",
  1172 => x"3f",
  1173 => x"20",
  1174 => x"24",
  1175 => x"6e",
  1176 => x"00",
  1177 => x"08",
  1178 => x"2a",
  1179 => x"2e",
  1180 => x"00",
  1181 => x"0c",
  1182 => x"20",
  1183 => x"2e",
  1184 => x"00",
  1185 => x"10",
  1186 => x"3e",
  1187 => x"00",
  1188 => x"76",
  1189 => x"00",
  1190 => x"36",
  1191 => x"00",
  1192 => x"28",
  1193 => x"05",
  1194 => x"42",
  1195 => x"44",
  1196 => x"88",
  1197 => x"83",
  1198 => x"48",
  1199 => x"43",
  1200 => x"42",
  1201 => x"43",
  1202 => x"86",
  1203 => x"45",
  1204 => x"24",
  1205 => x"85",
  1206 => x"34",
  1207 => x"80",
  1208 => x"24",
  1209 => x"12",
  1210 => x"b6",
  1211 => x"82",
  1212 => x"67",
  1213 => x"18",
  1214 => x"48",
  1215 => x"79",
  1216 => x"00",
  1217 => x"00",
  1218 => x"09",
  1219 => x"d2",
  1220 => x"4e",
  1221 => x"b9",
  1222 => x"00",
  1223 => x"00",
  1224 => x"03",
  1225 => x"0e",
  1226 => x"2f",
  1227 => x"02",
  1228 => x"4e",
  1229 => x"ba",
  1230 => x"fe",
  1231 => x"8e",
  1232 => x"b7",
  1233 => x"82",
  1234 => x"50",
  1235 => x"8f",
  1236 => x"60",
  1237 => x"02",
  1238 => x"74",
  1239 => x"00",
  1240 => x"2f",
  1241 => x"0a",
  1242 => x"4e",
  1243 => x"ba",
  1244 => x"fe",
  1245 => x"ea",
  1246 => x"2c",
  1247 => x"12",
  1248 => x"58",
  1249 => x"8f",
  1250 => x"b6",
  1251 => x"86",
  1252 => x"67",
  1253 => x"18",
  1254 => x"48",
  1255 => x"79",
  1256 => x"00",
  1257 => x"00",
  1258 => x"09",
  1259 => x"f6",
  1260 => x"4e",
  1261 => x"b9",
  1262 => x"00",
  1263 => x"00",
  1264 => x"03",
  1265 => x"0e",
  1266 => x"2f",
  1267 => x"06",
  1268 => x"4e",
  1269 => x"ba",
  1270 => x"fe",
  1271 => x"66",
  1272 => x"bd",
  1273 => x"83",
  1274 => x"84",
  1275 => x"83",
  1276 => x"50",
  1277 => x"8f",
  1278 => x"25",
  1279 => x"45",
  1280 => x"00",
  1281 => x"04",
  1282 => x"35",
  1283 => x"47",
  1284 => x"00",
  1285 => x"06",
  1286 => x"26",
  1287 => x"2a",
  1288 => x"00",
  1289 => x"04",
  1290 => x"b8",
  1291 => x"83",
  1292 => x"67",
  1293 => x"18",
  1294 => x"48",
  1295 => x"79",
  1296 => x"00",
  1297 => x"00",
  1298 => x"0a",
  1299 => x"1a",
  1300 => x"4e",
  1301 => x"b9",
  1302 => x"00",
  1303 => x"00",
  1304 => x"03",
  1305 => x"0e",
  1306 => x"2f",
  1307 => x"03",
  1308 => x"4e",
  1309 => x"ba",
  1310 => x"fe",
  1311 => x"3e",
  1312 => x"b9",
  1313 => x"83",
  1314 => x"84",
  1315 => x"83",
  1316 => x"50",
  1317 => x"8f",
  1318 => x"48",
  1319 => x"6a",
  1320 => x"00",
  1321 => x"04",
  1322 => x"4e",
  1323 => x"ba",
  1324 => x"fe",
  1325 => x"9a",
  1326 => x"26",
  1327 => x"2a",
  1328 => x"00",
  1329 => x"04",
  1330 => x"58",
  1331 => x"8f",
  1332 => x"b8",
  1333 => x"83",
  1334 => x"67",
  1335 => x"18",
  1336 => x"48",
  1337 => x"79",
  1338 => x"00",
  1339 => x"00",
  1340 => x"0a",
  1341 => x"3e",
  1342 => x"4e",
  1343 => x"b9",
  1344 => x"00",
  1345 => x"00",
  1346 => x"03",
  1347 => x"0e",
  1348 => x"2f",
  1349 => x"03",
  1350 => x"4e",
  1351 => x"ba",
  1352 => x"fe",
  1353 => x"14",
  1354 => x"b7",
  1355 => x"84",
  1356 => x"84",
  1357 => x"84",
  1358 => x"50",
  1359 => x"8f",
  1360 => x"20",
  1361 => x"02",
  1362 => x"4c",
  1363 => x"ee",
  1364 => x"04",
  1365 => x"fc",
  1366 => x"ff",
  1367 => x"e4",
  1368 => x"4e",
  1369 => x"5e",
  1370 => x"4e",
  1371 => x"75",
  1372 => x"4e",
  1373 => x"56",
  1374 => x"00",
  1375 => x"00",
  1376 => x"48",
  1377 => x"e7",
  1378 => x"3f",
  1379 => x"3c",
  1380 => x"24",
  1381 => x"6e",
  1382 => x"00",
  1383 => x"08",
  1384 => x"26",
  1385 => x"2e",
  1386 => x"00",
  1387 => x"0c",
  1388 => x"20",
  1389 => x"2e",
  1390 => x"00",
  1391 => x"10",
  1392 => x"78",
  1393 => x"00",
  1394 => x"18",
  1395 => x"00",
  1396 => x"72",
  1397 => x"ff",
  1398 => x"46",
  1399 => x"01",
  1400 => x"c2",
  1401 => x"83",
  1402 => x"82",
  1403 => x"84",
  1404 => x"28",
  1405 => x"41",
  1406 => x"2e",
  1407 => x"04",
  1408 => x"e1",
  1409 => x"8f",
  1410 => x"22",
  1411 => x"03",
  1412 => x"02",
  1413 => x"41",
  1414 => x"00",
  1415 => x"ff",
  1416 => x"8e",
  1417 => x"81",
  1418 => x"2c",
  1419 => x"04",
  1420 => x"48",
  1421 => x"46",
  1422 => x"42",
  1423 => x"46",
  1424 => x"22",
  1425 => x"03",
  1426 => x"02",
  1427 => x"81",
  1428 => x"ff",
  1429 => x"00",
  1430 => x"ff",
  1431 => x"ff",
  1432 => x"8c",
  1433 => x"81",
  1434 => x"2a",
  1435 => x"04",
  1436 => x"e1",
  1437 => x"4d",
  1438 => x"48",
  1439 => x"45",
  1440 => x"42",
  1441 => x"45",
  1442 => x"22",
  1443 => x"03",
  1444 => x"02",
  1445 => x"81",
  1446 => x"00",
  1447 => x"ff",
  1448 => x"ff",
  1449 => x"ff",
  1450 => x"8a",
  1451 => x"81",
  1452 => x"24",
  1453 => x"83",
  1454 => x"15",
  1455 => x"40",
  1456 => x"00",
  1457 => x"03",
  1458 => x"25",
  1459 => x"43",
  1460 => x"00",
  1461 => x"04",
  1462 => x"15",
  1463 => x"40",
  1464 => x"00",
  1465 => x"06",
  1466 => x"25",
  1467 => x"43",
  1468 => x"00",
  1469 => x"08",
  1470 => x"15",
  1471 => x"40",
  1472 => x"00",
  1473 => x"09",
  1474 => x"25",
  1475 => x"43",
  1476 => x"00",
  1477 => x"0c",
  1478 => x"15",
  1479 => x"40",
  1480 => x"00",
  1481 => x"0c",
  1482 => x"24",
  1483 => x"12",
  1484 => x"b9",
  1485 => x"c2",
  1486 => x"67",
  1487 => x"26",
  1488 => x"48",
  1489 => x"79",
  1490 => x"00",
  1491 => x"00",
  1492 => x"0a",
  1493 => x"62",
  1494 => x"4e",
  1495 => x"b9",
  1496 => x"00",
  1497 => x"00",
  1498 => x"03",
  1499 => x"0e",
  1500 => x"2f",
  1501 => x"02",
  1502 => x"47",
  1503 => x"fa",
  1504 => x"fd",
  1505 => x"7c",
  1506 => x"4e",
  1507 => x"93",
  1508 => x"2f",
  1509 => x"03",
  1510 => x"4e",
  1511 => x"93",
  1512 => x"2f",
  1513 => x"04",
  1514 => x"4e",
  1515 => x"93",
  1516 => x"20",
  1517 => x"0c",
  1518 => x"b1",
  1519 => x"82",
  1520 => x"4f",
  1521 => x"ef",
  1522 => x"00",
  1523 => x"10",
  1524 => x"60",
  1525 => x"02",
  1526 => x"74",
  1527 => x"00",
  1528 => x"47",
  1529 => x"ea",
  1530 => x"00",
  1531 => x"08",
  1532 => x"2f",
  1533 => x"0b",
  1534 => x"4e",
  1535 => x"ba",
  1536 => x"fd",
  1537 => x"c6",
  1538 => x"2a",
  1539 => x"52",
  1540 => x"58",
  1541 => x"8f",
  1542 => x"b9",
  1543 => x"cd",
  1544 => x"67",
  1545 => x"2a",
  1546 => x"48",
  1547 => x"79",
  1548 => x"00",
  1549 => x"00",
  1550 => x"0a",
  1551 => x"85",
  1552 => x"4e",
  1553 => x"b9",
  1554 => x"00",
  1555 => x"00",
  1556 => x"03",
  1557 => x"0e",
  1558 => x"2f",
  1559 => x"0d",
  1560 => x"4e",
  1561 => x"ba",
  1562 => x"fd",
  1563 => x"42",
  1564 => x"2f",
  1565 => x"03",
  1566 => x"4e",
  1567 => x"ba",
  1568 => x"fd",
  1569 => x"3c",
  1570 => x"2f",
  1571 => x"04",
  1572 => x"4e",
  1573 => x"ba",
  1574 => x"fd",
  1575 => x"36",
  1576 => x"20",
  1577 => x"0c",
  1578 => x"22",
  1579 => x"0d",
  1580 => x"b3",
  1581 => x"80",
  1582 => x"84",
  1583 => x"80",
  1584 => x"4f",
  1585 => x"ef",
  1586 => x"00",
  1587 => x"10",
  1588 => x"28",
  1589 => x"6a",
  1590 => x"00",
  1591 => x"04",
  1592 => x"be",
  1593 => x"8c",
  1594 => x"67",
  1595 => x"26",
  1596 => x"48",
  1597 => x"79",
  1598 => x"00",
  1599 => x"00",
  1600 => x"0a",
  1601 => x"a8",
  1602 => x"4e",
  1603 => x"b9",
  1604 => x"00",
  1605 => x"00",
  1606 => x"03",
  1607 => x"0e",
  1608 => x"2f",
  1609 => x"0c",
  1610 => x"4b",
  1611 => x"fa",
  1612 => x"fd",
  1613 => x"10",
  1614 => x"4e",
  1615 => x"95",
  1616 => x"2f",
  1617 => x"03",
  1618 => x"4e",
  1619 => x"95",
  1620 => x"2f",
  1621 => x"04",
  1622 => x"4e",
  1623 => x"95",
  1624 => x"20",
  1625 => x"0c",
  1626 => x"bf",
  1627 => x"80",
  1628 => x"84",
  1629 => x"80",
  1630 => x"4f",
  1631 => x"ef",
  1632 => x"00",
  1633 => x"10",
  1634 => x"2f",
  1635 => x"0b",
  1636 => x"4e",
  1637 => x"ba",
  1638 => x"fd",
  1639 => x"60",
  1640 => x"28",
  1641 => x"6a",
  1642 => x"00",
  1643 => x"04",
  1644 => x"58",
  1645 => x"8f",
  1646 => x"be",
  1647 => x"8c",
  1648 => x"67",
  1649 => x"26",
  1650 => x"48",
  1651 => x"79",
  1652 => x"00",
  1653 => x"00",
  1654 => x"0a",
  1655 => x"cb",
  1656 => x"4e",
  1657 => x"b9",
  1658 => x"00",
  1659 => x"00",
  1660 => x"03",
  1661 => x"0e",
  1662 => x"2f",
  1663 => x"0c",
  1664 => x"4b",
  1665 => x"fa",
  1666 => x"fc",
  1667 => x"da",
  1668 => x"4e",
  1669 => x"95",
  1670 => x"2f",
  1671 => x"03",
  1672 => x"4e",
  1673 => x"95",
  1674 => x"2f",
  1675 => x"04",
  1676 => x"4e",
  1677 => x"95",
  1678 => x"20",
  1679 => x"0c",
  1680 => x"b1",
  1681 => x"87",
  1682 => x"84",
  1683 => x"87",
  1684 => x"4f",
  1685 => x"ef",
  1686 => x"00",
  1687 => x"10",
  1688 => x"2e",
  1689 => x"2a",
  1690 => x"00",
  1691 => x"08",
  1692 => x"bc",
  1693 => x"87",
  1694 => x"67",
  1695 => x"24",
  1696 => x"48",
  1697 => x"79",
  1698 => x"00",
  1699 => x"00",
  1700 => x"0a",
  1701 => x"ee",
  1702 => x"4e",
  1703 => x"b9",
  1704 => x"00",
  1705 => x"00",
  1706 => x"03",
  1707 => x"0e",
  1708 => x"2f",
  1709 => x"07",
  1710 => x"49",
  1711 => x"fa",
  1712 => x"fc",
  1713 => x"ac",
  1714 => x"4e",
  1715 => x"94",
  1716 => x"2f",
  1717 => x"03",
  1718 => x"4e",
  1719 => x"94",
  1720 => x"2f",
  1721 => x"04",
  1722 => x"4e",
  1723 => x"94",
  1724 => x"bd",
  1725 => x"87",
  1726 => x"84",
  1727 => x"87",
  1728 => x"4f",
  1729 => x"ef",
  1730 => x"00",
  1731 => x"10",
  1732 => x"2f",
  1733 => x"0b",
  1734 => x"4e",
  1735 => x"ba",
  1736 => x"fc",
  1737 => x"fe",
  1738 => x"2e",
  1739 => x"2a",
  1740 => x"00",
  1741 => x"08",
  1742 => x"58",
  1743 => x"8f",
  1744 => x"bc",
  1745 => x"87",
  1746 => x"67",
  1747 => x"24",
  1748 => x"48",
  1749 => x"79",
  1750 => x"00",
  1751 => x"00",
  1752 => x"0b",
  1753 => x"11",
  1754 => x"4e",
  1755 => x"b9",
  1756 => x"00",
  1757 => x"00",
  1758 => x"03",
  1759 => x"0e",
  1760 => x"2f",
  1761 => x"07",
  1762 => x"49",
  1763 => x"fa",
  1764 => x"fc",
  1765 => x"78",
  1766 => x"4e",
  1767 => x"94",
  1768 => x"2f",
  1769 => x"03",
  1770 => x"4e",
  1771 => x"94",
  1772 => x"2f",
  1773 => x"04",
  1774 => x"4e",
  1775 => x"94",
  1776 => x"bf",
  1777 => x"86",
  1778 => x"84",
  1779 => x"86",
  1780 => x"4f",
  1781 => x"ef",
  1782 => x"00",
  1783 => x"10",
  1784 => x"2c",
  1785 => x"2a",
  1786 => x"00",
  1787 => x"0c",
  1788 => x"ba",
  1789 => x"86",
  1790 => x"67",
  1791 => x"24",
  1792 => x"48",
  1793 => x"79",
  1794 => x"00",
  1795 => x"00",
  1796 => x"0b",
  1797 => x"34",
  1798 => x"4e",
  1799 => x"b9",
  1800 => x"00",
  1801 => x"00",
  1802 => x"03",
  1803 => x"0e",
  1804 => x"2f",
  1805 => x"06",
  1806 => x"49",
  1807 => x"fa",
  1808 => x"fc",
  1809 => x"4c",
  1810 => x"4e",
  1811 => x"94",
  1812 => x"2f",
  1813 => x"03",
  1814 => x"4e",
  1815 => x"94",
  1816 => x"2f",
  1817 => x"04",
  1818 => x"4e",
  1819 => x"94",
  1820 => x"bb",
  1821 => x"86",
  1822 => x"84",
  1823 => x"86",
  1824 => x"4f",
  1825 => x"ef",
  1826 => x"00",
  1827 => x"10",
  1828 => x"2f",
  1829 => x"0b",
  1830 => x"4e",
  1831 => x"ba",
  1832 => x"fc",
  1833 => x"9e",
  1834 => x"2c",
  1835 => x"2a",
  1836 => x"00",
  1837 => x"0c",
  1838 => x"58",
  1839 => x"8f",
  1840 => x"ba",
  1841 => x"86",
  1842 => x"67",
  1843 => x"24",
  1844 => x"48",
  1845 => x"79",
  1846 => x"00",
  1847 => x"00",
  1848 => x"0b",
  1849 => x"57",
  1850 => x"4e",
  1851 => x"b9",
  1852 => x"00",
  1853 => x"00",
  1854 => x"03",
  1855 => x"0e",
  1856 => x"2f",
  1857 => x"06",
  1858 => x"45",
  1859 => x"fa",
  1860 => x"fc",
  1861 => x"18",
  1862 => x"4e",
  1863 => x"92",
  1864 => x"2f",
  1865 => x"03",
  1866 => x"4e",
  1867 => x"92",
  1868 => x"2f",
  1869 => x"04",
  1870 => x"4e",
  1871 => x"92",
  1872 => x"bd",
  1873 => x"85",
  1874 => x"84",
  1875 => x"85",
  1876 => x"4f",
  1877 => x"ef",
  1878 => x"00",
  1879 => x"10",
  1880 => x"20",
  1881 => x"02",
  1882 => x"4c",
  1883 => x"ee",
  1884 => x"3c",
  1885 => x"fc",
  1886 => x"ff",
  1887 => x"d8",
  1888 => x"4e",
  1889 => x"5e",
  1890 => x"4e",
  1891 => x"75",
  1892 => x"4e",
  1893 => x"56",
  1894 => x"00",
  1895 => x"00",
  1896 => x"48",
  1897 => x"e7",
  1898 => x"3f",
  1899 => x"30",
  1900 => x"2e",
  1901 => x"2e",
  1902 => x"00",
  1903 => x"08",
  1904 => x"48",
  1905 => x"79",
  1906 => x"00",
  1907 => x"00",
  1908 => x"0b",
  1909 => x"7a",
  1910 => x"4e",
  1911 => x"b9",
  1912 => x"00",
  1913 => x"00",
  1914 => x"03",
  1915 => x"0e",
  1916 => x"58",
  1917 => x"8f",
  1918 => x"76",
  1919 => x"00",
  1920 => x"74",
  1921 => x"00",
  1922 => x"47",
  1923 => x"fa",
  1924 => x"fd",
  1925 => x"0a",
  1926 => x"45",
  1927 => x"f9",
  1928 => x"00",
  1929 => x"00",
  1930 => x"02",
  1931 => x"f0",
  1932 => x"60",
  1933 => x"34",
  1934 => x"3f",
  1935 => x"04",
  1936 => x"42",
  1937 => x"67",
  1938 => x"2f",
  1939 => x"03",
  1940 => x"2f",
  1941 => x"07",
  1942 => x"4e",
  1943 => x"93",
  1944 => x"84",
  1945 => x"80",
  1946 => x"06",
  1947 => x"84",
  1948 => x"00",
  1949 => x"31",
  1950 => x"87",
  1951 => x"65",
  1952 => x"4f",
  1953 => x"ef",
  1954 => x"00",
  1955 => x"0c",
  1956 => x"0c",
  1957 => x"84",
  1958 => x"80",
  1959 => x"14",
  1960 => x"1f",
  1961 => x"2e",
  1962 => x"66",
  1963 => x"e2",
  1964 => x"48",
  1965 => x"78",
  1966 => x"00",
  1967 => x"2e",
  1968 => x"4e",
  1969 => x"92",
  1970 => x"06",
  1971 => x"83",
  1972 => x"00",
  1973 => x"21",
  1974 => x"23",
  1975 => x"45",
  1976 => x"58",
  1977 => x"8f",
  1978 => x"0c",
  1979 => x"83",
  1980 => x"80",
  1981 => x"05",
  1982 => x"41",
  1983 => x"91",
  1984 => x"67",
  1985 => x"04",
  1986 => x"78",
  1987 => x"00",
  1988 => x"60",
  1989 => x"c8",
  1990 => x"4a",
  1991 => x"82",
  1992 => x"67",
  1993 => x"18",
  1994 => x"48",
  1995 => x"79",
  1996 => x"00",
  1997 => x"00",
  1998 => x"0b",
  1999 => x"8f",
  2000 => x"4e",
  2001 => x"b9",
  2002 => x"00",
  2003 => x"00",
  2004 => x"03",
  2005 => x"0e",
  2006 => x"2f",
  2007 => x"02",
  2008 => x"4e",
  2009 => x"ba",
  2010 => x"fb",
  2011 => x"82",
  2012 => x"50",
  2013 => x"8f",
  2014 => x"78",
  2015 => x"00",
  2016 => x"60",
  2017 => x"02",
  2018 => x"78",
  2019 => x"01",
  2020 => x"48",
  2021 => x"79",
  2022 => x"00",
  2023 => x"00",
  2024 => x"0b",
  2025 => x"af",
  2026 => x"4e",
  2027 => x"b9",
  2028 => x"00",
  2029 => x"00",
  2030 => x"03",
  2031 => x"0e",
  2032 => x"58",
  2033 => x"8f",
  2034 => x"7a",
  2035 => x"00",
  2036 => x"76",
  2037 => x"00",
  2038 => x"47",
  2039 => x"fa",
  2040 => x"fc",
  2041 => x"1c",
  2042 => x"45",
  2043 => x"f9",
  2044 => x"00",
  2045 => x"00",
  2046 => x"02",
  2047 => x"f0",
  2048 => x"60",
  2049 => x"32",
  2050 => x"2f",
  2051 => x"06",
  2052 => x"2f",
  2053 => x"05",
  2054 => x"2f",
  2055 => x"07",
  2056 => x"4e",
  2057 => x"93",
  2058 => x"86",
  2059 => x"80",
  2060 => x"06",
  2061 => x"86",
  2062 => x"00",
  2063 => x"19",
  2064 => x"87",
  2065 => x"65",
  2066 => x"4f",
  2067 => x"ef",
  2068 => x"00",
  2069 => x"0c",
  2070 => x"0c",
  2071 => x"86",
  2072 => x"80",
  2073 => x"0b",
  2074 => x"16",
  2075 => x"94",
  2076 => x"66",
  2077 => x"e4",
  2078 => x"48",
  2079 => x"78",
  2080 => x"00",
  2081 => x"2e",
  2082 => x"4e",
  2083 => x"92",
  2084 => x"06",
  2085 => x"85",
  2086 => x"00",
  2087 => x"13",
  2088 => x"45",
  2089 => x"67",
  2090 => x"58",
  2091 => x"8f",
  2092 => x"0c",
  2093 => x"85",
  2094 => x"80",
  2095 => x"0c",
  2096 => x"25",
  2097 => x"63",
  2098 => x"67",
  2099 => x"04",
  2100 => x"7c",
  2101 => x"00",
  2102 => x"60",
  2103 => x"ca",
  2104 => x"4a",
  2105 => x"83",
  2106 => x"67",
  2107 => x"0a",
  2108 => x"2f",
  2109 => x"03",
  2110 => x"4e",
  2111 => x"ba",
  2112 => x"fb",
  2113 => x"1c",
  2114 => x"58",
  2115 => x"8f",
  2116 => x"78",
  2117 => x"00",
  2118 => x"86",
  2119 => x"82",
  2120 => x"48",
  2121 => x"79",
  2122 => x"00",
  2123 => x"00",
  2124 => x"0b",
  2125 => x"c9",
  2126 => x"4e",
  2127 => x"b9",
  2128 => x"00",
  2129 => x"00",
  2130 => x"03",
  2131 => x"0e",
  2132 => x"58",
  2133 => x"8f",
  2134 => x"7a",
  2135 => x"00",
  2136 => x"74",
  2137 => x"00",
  2138 => x"47",
  2139 => x"fa",
  2140 => x"fd",
  2141 => x"00",
  2142 => x"45",
  2143 => x"f9",
  2144 => x"00",
  2145 => x"00",
  2146 => x"02",
  2147 => x"f0",
  2148 => x"60",
  2149 => x"36",
  2150 => x"70",
  2151 => x"00",
  2152 => x"10",
  2153 => x"06",
  2154 => x"2f",
  2155 => x"00",
  2156 => x"2f",
  2157 => x"05",
  2158 => x"2f",
  2159 => x"07",
  2160 => x"4e",
  2161 => x"93",
  2162 => x"84",
  2163 => x"80",
  2164 => x"06",
  2165 => x"86",
  2166 => x"00",
  2167 => x"28",
  2168 => x"76",
  2169 => x"53",
  2170 => x"4f",
  2171 => x"ef",
  2172 => x"00",
  2173 => x"0c",
  2174 => x"0c",
  2175 => x"86",
  2176 => x"80",
  2177 => x"06",
  2178 => x"62",
  2179 => x"9e",
  2180 => x"66",
  2181 => x"e0",
  2182 => x"48",
  2183 => x"78",
  2184 => x"00",
  2185 => x"2e",
  2186 => x"4e",
  2187 => x"92",
  2188 => x"06",
  2189 => x"85",
  2190 => x"00",
  2191 => x"71",
  2192 => x"23",
  2193 => x"41",
  2194 => x"58",
  2195 => x"8f",
  2196 => x"0c",
  2197 => x"85",
  2198 => x"80",
  2199 => x"29",
  2200 => x"ef",
  2201 => x"a2",
  2202 => x"67",
  2203 => x"04",
  2204 => x"7c",
  2205 => x"00",
  2206 => x"60",
  2207 => x"c6",
  2208 => x"4a",
  2209 => x"82",
  2210 => x"67",
  2211 => x"0a",
  2212 => x"2f",
  2213 => x"02",
  2214 => x"4e",
  2215 => x"ba",
  2216 => x"fa",
  2217 => x"b4",
  2218 => x"58",
  2219 => x"8f",
  2220 => x"78",
  2221 => x"00",
  2222 => x"84",
  2223 => x"83",
  2224 => x"67",
  2225 => x"14",
  2226 => x"48",
  2227 => x"79",
  2228 => x"00",
  2229 => x"00",
  2230 => x"0b",
  2231 => x"de",
  2232 => x"4e",
  2233 => x"b9",
  2234 => x"00",
  2235 => x"00",
  2236 => x"03",
  2237 => x"0e",
  2238 => x"2f",
  2239 => x"02",
  2240 => x"4e",
  2241 => x"ba",
  2242 => x"fa",
  2243 => x"9a",
  2244 => x"50",
  2245 => x"8f",
  2246 => x"20",
  2247 => x"04",
  2248 => x"4c",
  2249 => x"ee",
  2250 => x"0c",
  2251 => x"fc",
  2252 => x"ff",
  2253 => x"e0",
  2254 => x"4e",
  2255 => x"5e",
  2256 => x"4e",
  2257 => x"75",
  2258 => x"00",
  2259 => x"00",
  2260 => x"30",
  2261 => x"2f",
  2262 => x"00",
  2263 => x"04",
  2264 => x"c0",
  2265 => x"ef",
  2266 => x"00",
  2267 => x"0a",
  2268 => x"32",
  2269 => x"2f",
  2270 => x"00",
  2271 => x"06",
  2272 => x"c2",
  2273 => x"ef",
  2274 => x"00",
  2275 => x"08",
  2276 => x"d0",
  2277 => x"41",
  2278 => x"48",
  2279 => x"40",
  2280 => x"42",
  2281 => x"40",
  2282 => x"32",
  2283 => x"2f",
  2284 => x"00",
  2285 => x"06",
  2286 => x"c2",
  2287 => x"ef",
  2288 => x"00",
  2289 => x"0a",
  2290 => x"d0",
  2291 => x"81",
  2292 => x"4e",
  2293 => x"75",
  2294 => x"00",
  2295 => x"00",
  2296 => x"2f",
  2297 => x"02",
  2298 => x"74",
  2299 => x"01",
  2300 => x"22",
  2301 => x"2f",
  2302 => x"00",
  2303 => x"0c",
  2304 => x"6a",
  2305 => x"04",
  2306 => x"44",
  2307 => x"81",
  2308 => x"44",
  2309 => x"02",
  2310 => x"20",
  2311 => x"2f",
  2312 => x"00",
  2313 => x"08",
  2314 => x"6a",
  2315 => x"04",
  2316 => x"44",
  2317 => x"80",
  2318 => x"44",
  2319 => x"02",
  2320 => x"2f",
  2321 => x"01",
  2322 => x"2f",
  2323 => x"00",
  2324 => x"4e",
  2325 => x"b9",
  2326 => x"00",
  2327 => x"00",
  2328 => x"09",
  2329 => x"28",
  2330 => x"50",
  2331 => x"8f",
  2332 => x"4a",
  2333 => x"02",
  2334 => x"6a",
  2335 => x"02",
  2336 => x"44",
  2337 => x"80",
  2338 => x"24",
  2339 => x"1f",
  2340 => x"4e",
  2341 => x"75",
  2342 => x"00",
  2343 => x"00",
  2344 => x"2f",
  2345 => x"02",
  2346 => x"22",
  2347 => x"2f",
  2348 => x"00",
  2349 => x"0c",
  2350 => x"20",
  2351 => x"2f",
  2352 => x"00",
  2353 => x"08",
  2354 => x"0c",
  2355 => x"81",
  2356 => x"00",
  2357 => x"01",
  2358 => x"00",
  2359 => x"00",
  2360 => x"64",
  2361 => x"16",
  2362 => x"24",
  2363 => x"00",
  2364 => x"42",
  2365 => x"42",
  2366 => x"48",
  2367 => x"42",
  2368 => x"84",
  2369 => x"c1",
  2370 => x"30",
  2371 => x"02",
  2372 => x"48",
  2373 => x"40",
  2374 => x"34",
  2375 => x"2f",
  2376 => x"00",
  2377 => x"0a",
  2378 => x"84",
  2379 => x"c1",
  2380 => x"30",
  2381 => x"02",
  2382 => x"60",
  2383 => x"30",
  2384 => x"24",
  2385 => x"01",
  2386 => x"e2",
  2387 => x"89",
  2388 => x"e2",
  2389 => x"88",
  2390 => x"0c",
  2391 => x"81",
  2392 => x"00",
  2393 => x"01",
  2394 => x"00",
  2395 => x"00",
  2396 => x"64",
  2397 => x"f4",
  2398 => x"80",
  2399 => x"c1",
  2400 => x"02",
  2401 => x"80",
  2402 => x"00",
  2403 => x"00",
  2404 => x"ff",
  2405 => x"ff",
  2406 => x"22",
  2407 => x"02",
  2408 => x"c2",
  2409 => x"c0",
  2410 => x"48",
  2411 => x"42",
  2412 => x"c4",
  2413 => x"c0",
  2414 => x"48",
  2415 => x"42",
  2416 => x"4a",
  2417 => x"42",
  2418 => x"66",
  2419 => x"0a",
  2420 => x"d2",
  2421 => x"82",
  2422 => x"65",
  2423 => x"06",
  2424 => x"b2",
  2425 => x"af",
  2426 => x"00",
  2427 => x"08",
  2428 => x"63",
  2429 => x"02",
  2430 => x"53",
  2431 => x"80",
  2432 => x"24",
  2433 => x"1f",
  2434 => x"4e",
  2435 => x"75",
  2436 => x"4d",
  2437 => x"69",
  2438 => x"73",
  2439 => x"61",
  2440 => x"6c",
  2441 => x"69",
  2442 => x"67",
  2443 => x"6e",
  2444 => x"65",
  2445 => x"64",
  2446 => x"20",
  2447 => x"6c",
  2448 => x"6f",
  2449 => x"6e",
  2450 => x"67",
  2451 => x"20",
  2452 => x"63",
  2453 => x"68",
  2454 => x"65",
  2455 => x"63",
  2456 => x"6b",
  2457 => x"20",
  2458 => x"28",
  2459 => x"63",
  2460 => x"61",
  2461 => x"63",
  2462 => x"68",
  2463 => x"65",
  2464 => x"29",
  2465 => x"20",
  2466 => x"66",
  2467 => x"61",
  2468 => x"69",
  2469 => x"6c",
  2470 => x"65",
  2471 => x"64",
  2472 => x"3a",
  2473 => x"20",
  2474 => x"00",
  2475 => x"4d",
  2476 => x"69",
  2477 => x"73",
  2478 => x"61",
  2479 => x"6c",
  2480 => x"69",
  2481 => x"67",
  2482 => x"6e",
  2483 => x"65",
  2484 => x"64",
  2485 => x"20",
  2486 => x"6c",
  2487 => x"6f",
  2488 => x"6e",
  2489 => x"67",
  2490 => x"20",
  2491 => x"63",
  2492 => x"68",
  2493 => x"65",
  2494 => x"63",
  2495 => x"6b",
  2496 => x"20",
  2497 => x"28",
  2498 => x"66",
  2499 => x"6c",
  2500 => x"75",
  2501 => x"73",
  2502 => x"68",
  2503 => x"29",
  2504 => x"20",
  2505 => x"66",
  2506 => x"61",
  2507 => x"69",
  2508 => x"6c",
  2509 => x"65",
  2510 => x"64",
  2511 => x"3a",
  2512 => x"20",
  2513 => x"00",
  2514 => x"4c",
  2515 => x"6f",
  2516 => x"6e",
  2517 => x"67",
  2518 => x"20",
  2519 => x"53",
  2520 => x"68",
  2521 => x"6f",
  2522 => x"72",
  2523 => x"74",
  2524 => x"20",
  2525 => x"63",
  2526 => x"68",
  2527 => x"65",
  2528 => x"63",
  2529 => x"6b",
  2530 => x"20",
  2531 => x"31",
  2532 => x"20",
  2533 => x"28",
  2534 => x"63",
  2535 => x"61",
  2536 => x"63",
  2537 => x"68",
  2538 => x"65",
  2539 => x"29",
  2540 => x"20",
  2541 => x"66",
  2542 => x"61",
  2543 => x"69",
  2544 => x"6c",
  2545 => x"65",
  2546 => x"64",
  2547 => x"3a",
  2548 => x"20",
  2549 => x"00",
  2550 => x"4c",
  2551 => x"6f",
  2552 => x"6e",
  2553 => x"67",
  2554 => x"20",
  2555 => x"53",
  2556 => x"68",
  2557 => x"6f",
  2558 => x"72",
  2559 => x"74",
  2560 => x"20",
  2561 => x"63",
  2562 => x"68",
  2563 => x"65",
  2564 => x"63",
  2565 => x"6b",
  2566 => x"20",
  2567 => x"31",
  2568 => x"20",
  2569 => x"28",
  2570 => x"66",
  2571 => x"6c",
  2572 => x"75",
  2573 => x"73",
  2574 => x"68",
  2575 => x"29",
  2576 => x"20",
  2577 => x"66",
  2578 => x"61",
  2579 => x"69",
  2580 => x"6c",
  2581 => x"65",
  2582 => x"64",
  2583 => x"3a",
  2584 => x"20",
  2585 => x"00",
  2586 => x"4c",
  2587 => x"6f",
  2588 => x"6e",
  2589 => x"67",
  2590 => x"20",
  2591 => x"53",
  2592 => x"68",
  2593 => x"6f",
  2594 => x"72",
  2595 => x"74",
  2596 => x"20",
  2597 => x"63",
  2598 => x"68",
  2599 => x"65",
  2600 => x"63",
  2601 => x"6b",
  2602 => x"20",
  2603 => x"32",
  2604 => x"20",
  2605 => x"28",
  2606 => x"63",
  2607 => x"61",
  2608 => x"63",
  2609 => x"68",
  2610 => x"65",
  2611 => x"29",
  2612 => x"20",
  2613 => x"66",
  2614 => x"61",
  2615 => x"69",
  2616 => x"6c",
  2617 => x"65",
  2618 => x"64",
  2619 => x"3a",
  2620 => x"20",
  2621 => x"00",
  2622 => x"4c",
  2623 => x"6f",
  2624 => x"6e",
  2625 => x"67",
  2626 => x"20",
  2627 => x"53",
  2628 => x"68",
  2629 => x"6f",
  2630 => x"72",
  2631 => x"74",
  2632 => x"20",
  2633 => x"63",
  2634 => x"68",
  2635 => x"65",
  2636 => x"63",
  2637 => x"6b",
  2638 => x"20",
  2639 => x"32",
  2640 => x"20",
  2641 => x"28",
  2642 => x"66",
  2643 => x"6c",
  2644 => x"75",
  2645 => x"73",
  2646 => x"68",
  2647 => x"29",
  2648 => x"20",
  2649 => x"66",
  2650 => x"61",
  2651 => x"69",
  2652 => x"6c",
  2653 => x"65",
  2654 => x"64",
  2655 => x"3a",
  2656 => x"20",
  2657 => x"00",
  2658 => x"4c",
  2659 => x"6f",
  2660 => x"6e",
  2661 => x"67",
  2662 => x"20",
  2663 => x"42",
  2664 => x"79",
  2665 => x"74",
  2666 => x"65",
  2667 => x"20",
  2668 => x"63",
  2669 => x"68",
  2670 => x"65",
  2671 => x"63",
  2672 => x"6b",
  2673 => x"20",
  2674 => x"31",
  2675 => x"20",
  2676 => x"28",
  2677 => x"63",
  2678 => x"61",
  2679 => x"63",
  2680 => x"68",
  2681 => x"65",
  2682 => x"29",
  2683 => x"20",
  2684 => x"66",
  2685 => x"61",
  2686 => x"69",
  2687 => x"6c",
  2688 => x"65",
  2689 => x"64",
  2690 => x"3a",
  2691 => x"20",
  2692 => x"00",
  2693 => x"4c",
  2694 => x"6f",
  2695 => x"6e",
  2696 => x"67",
  2697 => x"20",
  2698 => x"42",
  2699 => x"79",
  2700 => x"74",
  2701 => x"65",
  2702 => x"20",
  2703 => x"63",
  2704 => x"68",
  2705 => x"65",
  2706 => x"63",
  2707 => x"6b",
  2708 => x"20",
  2709 => x"31",
  2710 => x"20",
  2711 => x"28",
  2712 => x"66",
  2713 => x"6c",
  2714 => x"75",
  2715 => x"73",
  2716 => x"68",
  2717 => x"29",
  2718 => x"20",
  2719 => x"66",
  2720 => x"61",
  2721 => x"69",
  2722 => x"6c",
  2723 => x"65",
  2724 => x"64",
  2725 => x"3a",
  2726 => x"20",
  2727 => x"00",
  2728 => x"4c",
  2729 => x"6f",
  2730 => x"6e",
  2731 => x"67",
  2732 => x"20",
  2733 => x"42",
  2734 => x"79",
  2735 => x"74",
  2736 => x"65",
  2737 => x"20",
  2738 => x"63",
  2739 => x"68",
  2740 => x"65",
  2741 => x"63",
  2742 => x"6b",
  2743 => x"20",
  2744 => x"32",
  2745 => x"20",
  2746 => x"28",
  2747 => x"63",
  2748 => x"61",
  2749 => x"63",
  2750 => x"68",
  2751 => x"65",
  2752 => x"29",
  2753 => x"20",
  2754 => x"66",
  2755 => x"61",
  2756 => x"69",
  2757 => x"6c",
  2758 => x"65",
  2759 => x"64",
  2760 => x"3a",
  2761 => x"20",
  2762 => x"00",
  2763 => x"4c",
  2764 => x"6f",
  2765 => x"6e",
  2766 => x"67",
  2767 => x"20",
  2768 => x"42",
  2769 => x"79",
  2770 => x"74",
  2771 => x"65",
  2772 => x"20",
  2773 => x"63",
  2774 => x"68",
  2775 => x"65",
  2776 => x"63",
  2777 => x"6b",
  2778 => x"20",
  2779 => x"32",
  2780 => x"20",
  2781 => x"28",
  2782 => x"66",
  2783 => x"6c",
  2784 => x"75",
  2785 => x"73",
  2786 => x"68",
  2787 => x"29",
  2788 => x"20",
  2789 => x"66",
  2790 => x"61",
  2791 => x"69",
  2792 => x"6c",
  2793 => x"65",
  2794 => x"64",
  2795 => x"3a",
  2796 => x"20",
  2797 => x"00",
  2798 => x"4c",
  2799 => x"6f",
  2800 => x"6e",
  2801 => x"67",
  2802 => x"20",
  2803 => x"42",
  2804 => x"79",
  2805 => x"74",
  2806 => x"65",
  2807 => x"20",
  2808 => x"63",
  2809 => x"68",
  2810 => x"65",
  2811 => x"63",
  2812 => x"6b",
  2813 => x"20",
  2814 => x"33",
  2815 => x"20",
  2816 => x"28",
  2817 => x"63",
  2818 => x"61",
  2819 => x"63",
  2820 => x"68",
  2821 => x"65",
  2822 => x"29",
  2823 => x"20",
  2824 => x"66",
  2825 => x"61",
  2826 => x"69",
  2827 => x"6c",
  2828 => x"65",
  2829 => x"64",
  2830 => x"3a",
  2831 => x"20",
  2832 => x"00",
  2833 => x"4c",
  2834 => x"6f",
  2835 => x"6e",
  2836 => x"67",
  2837 => x"20",
  2838 => x"42",
  2839 => x"79",
  2840 => x"74",
  2841 => x"65",
  2842 => x"20",
  2843 => x"63",
  2844 => x"68",
  2845 => x"65",
  2846 => x"63",
  2847 => x"6b",
  2848 => x"20",
  2849 => x"33",
  2850 => x"20",
  2851 => x"28",
  2852 => x"66",
  2853 => x"6c",
  2854 => x"75",
  2855 => x"73",
  2856 => x"68",
  2857 => x"29",
  2858 => x"20",
  2859 => x"66",
  2860 => x"61",
  2861 => x"69",
  2862 => x"6c",
  2863 => x"65",
  2864 => x"64",
  2865 => x"3a",
  2866 => x"20",
  2867 => x"00",
  2868 => x"4c",
  2869 => x"6f",
  2870 => x"6e",
  2871 => x"67",
  2872 => x"20",
  2873 => x"42",
  2874 => x"79",
  2875 => x"74",
  2876 => x"65",
  2877 => x"20",
  2878 => x"63",
  2879 => x"68",
  2880 => x"65",
  2881 => x"63",
  2882 => x"6b",
  2883 => x"20",
  2884 => x"34",
  2885 => x"20",
  2886 => x"28",
  2887 => x"63",
  2888 => x"61",
  2889 => x"63",
  2890 => x"68",
  2891 => x"65",
  2892 => x"29",
  2893 => x"20",
  2894 => x"66",
  2895 => x"61",
  2896 => x"69",
  2897 => x"6c",
  2898 => x"65",
  2899 => x"64",
  2900 => x"3a",
  2901 => x"20",
  2902 => x"00",
  2903 => x"4c",
  2904 => x"6f",
  2905 => x"6e",
  2906 => x"67",
  2907 => x"20",
  2908 => x"42",
  2909 => x"79",
  2910 => x"74",
  2911 => x"65",
  2912 => x"20",
  2913 => x"63",
  2914 => x"68",
  2915 => x"65",
  2916 => x"63",
  2917 => x"6b",
  2918 => x"20",
  2919 => x"34",
  2920 => x"20",
  2921 => x"28",
  2922 => x"66",
  2923 => x"6c",
  2924 => x"75",
  2925 => x"73",
  2926 => x"68",
  2927 => x"29",
  2928 => x"20",
  2929 => x"66",
  2930 => x"61",
  2931 => x"69",
  2932 => x"6c",
  2933 => x"65",
  2934 => x"64",
  2935 => x"3a",
  2936 => x"20",
  2937 => x"00",
  2938 => x"0a",
  2939 => x"4c",
  2940 => x"6f",
  2941 => x"6e",
  2942 => x"67",
  2943 => x"2f",
  2944 => x"73",
  2945 => x"68",
  2946 => x"6f",
  2947 => x"72",
  2948 => x"74",
  2949 => x"20",
  2950 => x"74",
  2951 => x"65",
  2952 => x"73",
  2953 => x"74",
  2954 => x"2e",
  2955 => x"2e",
  2956 => x"2e",
  2957 => x"0a",
  2958 => x"00",
  2959 => x"42",
  2960 => x"61",
  2961 => x"64",
  2962 => x"20",
  2963 => x"62",
  2964 => x"69",
  2965 => x"74",
  2966 => x"73",
  2967 => x"20",
  2968 => x"66",
  2969 => x"72",
  2970 => x"6f",
  2971 => x"6d",
  2972 => x"20",
  2973 => x"4c",
  2974 => x"6f",
  2975 => x"6e",
  2976 => x"67",
  2977 => x"20",
  2978 => x"53",
  2979 => x"68",
  2980 => x"6f",
  2981 => x"72",
  2982 => x"74",
  2983 => x"20",
  2984 => x"74",
  2985 => x"65",
  2986 => x"73",
  2987 => x"74",
  2988 => x"3a",
  2989 => x"20",
  2990 => x"00",
  2991 => x"0a",
  2992 => x"4d",
  2993 => x"69",
  2994 => x"73",
  2995 => x"61",
  2996 => x"6c",
  2997 => x"69",
  2998 => x"67",
  2999 => x"6e",
  3000 => x"65",
  3001 => x"64",
  3002 => x"20",
  3003 => x"4c",
  3004 => x"6f",
  3005 => x"6e",
  3006 => x"67",
  3007 => x"20",
  3008 => x"74",
  3009 => x"65",
  3010 => x"73",
  3011 => x"74",
  3012 => x"2e",
  3013 => x"2e",
  3014 => x"2e",
  3015 => x"0a",
  3016 => x"00",
  3017 => x"4c",
  3018 => x"6f",
  3019 => x"6e",
  3020 => x"67",
  3021 => x"20",
  3022 => x"2f",
  3023 => x"20",
  3024 => x"62",
  3025 => x"79",
  3026 => x"74",
  3027 => x"65",
  3028 => x"20",
  3029 => x"74",
  3030 => x"65",
  3031 => x"73",
  3032 => x"74",
  3033 => x"2e",
  3034 => x"2e",
  3035 => x"2e",
  3036 => x"0a",
  3037 => x"00",
  3038 => x"42",
  3039 => x"61",
  3040 => x"64",
  3041 => x"20",
  3042 => x"62",
  3043 => x"69",
  3044 => x"74",
  3045 => x"73",
  3046 => x"20",
  3047 => x"64",
  3048 => x"65",
  3049 => x"74",
  3050 => x"65",
  3051 => x"63",
  3052 => x"74",
  3053 => x"65",
  3054 => x"64",
  3055 => x"3a",
  3056 => x"20",
  3057 => x"00",
  3058 => x"48",
  3059 => x"65",
  3060 => x"6c",
  3061 => x"6c",
  3062 => x"6f",
  3063 => x"2c",
  3064 => x"20",
  3065 => x"77",
  3066 => x"6f",
  3067 => x"72",
  3068 => x"6c",
  3069 => x"64",
  3070 => x"21",
  3071 => x"00",
  3072 => x"43",
  3073 => x"6f",
  3074 => x"6d",
  3075 => x"6d",
  3076 => x"65",
  3077 => x"6e",
  3078 => x"63",
  3079 => x"69",
  3080 => x"6e",
  3081 => x"67",
  3082 => x"20",
  3083 => x"73",
  3084 => x"61",
  3085 => x"6e",
  3086 => x"69",
  3087 => x"74",
  3088 => x"79",
  3089 => x"20",
  3090 => x"63",
  3091 => x"68",
  3092 => x"65",
  3093 => x"63",
  3094 => x"6b",
  3095 => x"73",
  3096 => x"2e",
  3097 => x"2e",
  3098 => x"2e",
  3099 => x"0a",
  3100 => x"00",
  3101 => x"4d",
  3102 => x"65",
  3103 => x"6d",
  3104 => x"6f",
  3105 => x"72",
  3106 => x"79",
  3107 => x"20",
  3108 => x"63",
  3109 => x"68",
  3110 => x"65",
  3111 => x"63",
  3112 => x"6b",
  3113 => x"20",
  3114 => x"70",
  3115 => x"61",
  3116 => x"73",
  3117 => x"73",
  3118 => x"65",
  3119 => x"64",
  3120 => x"0a",
  3121 => x"00",
  3122 => x"4d",
  3123 => x"65",
  3124 => x"6d",
  3125 => x"6f",
  3126 => x"72",
  3127 => x"79",
  3128 => x"20",
  3129 => x"63",
  3130 => x"68",
  3131 => x"65",
  3132 => x"63",
  3133 => x"6b",
  3134 => x"20",
  3135 => x"66",
  3136 => x"61",
  3137 => x"69",
  3138 => x"6c",
  3139 => x"65",
  3140 => x"64",
  3141 => x"0a",
  3142 => x"00",
  3143 => x"00",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

